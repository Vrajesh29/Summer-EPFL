module adderTree2(
  input         clock,
  input         reset,
  input  [5:0]  io_sign_man_0,
  input  [5:0]  io_sign_man_1,
  input  [5:0]  io_sign_man_2,
  input  [5:0]  io_sign_man_3,
  input  [8:0]  io_exps_0,
  input  [8:0]  io_exps_1,
  input  [8:0]  io_exps_2,
  input  [8:0]  io_exps_3,
  input         io_control_signal,
  input         io_control_signal2,
  output [13:0] io_result_tree
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] exp_buffer_0; // @[block_division.scala 243:60]
  reg [8:0] exp_buffer_1; // @[block_division.scala 243:60]
  reg [8:0] exp_buffer_2; // @[block_division.scala 243:60]
  reg [8:0] exp_buffer_3; // @[block_division.scala 243:60]
  reg [5:0] man_buffer_two_complement_0; // @[block_division.scala 245:12]
  reg [5:0] man_buffer_two_complement_1; // @[block_division.scala 245:12]
  reg [5:0] man_buffer_two_complement_2; // @[block_division.scala 245:12]
  reg [5:0] man_buffer_two_complement_3; // @[block_division.scala 245:12]
  wire [5:0] _GEN_1 = ~io_control_signal ? $signed(io_sign_man_0) : $signed(man_buffer_two_complement_0); // @[block_division.scala 245:12 249:34 253:36]
  wire [5:0] _GEN_3 = ~io_control_signal ? $signed(io_sign_man_1) : $signed(man_buffer_two_complement_1); // @[block_division.scala 245:12 249:34 253:36]
  reg [9:0] v; // @[block_division.scala 259:18]
  reg  enable; // @[block_division.scala 260:19]
  wire  _GEN_8 = io_control_signal2 | enable; // @[block_division.scala 261:36 262:12 260:19]
  wire [9:0] _v_T_1 = v + 10'h1; // @[block_division.scala 270:16]
  wire  _exp_buffer_0_T = exp_buffer_0 > exp_buffer_1; // @[block_division.scala 274:31]
  wire [8:0] _exp_difference_T_2 = exp_buffer_0 - exp_buffer_1; // @[block_division.scala 280:31]
  wire [8:0] _exp_difference_T_4 = exp_buffer_1 - exp_buffer_0; // @[block_division.scala 281:35]
  wire [8:0] exp_difference = _exp_buffer_0_T ? _exp_difference_T_2 : _exp_difference_T_4; // @[block_division.scala 278:35]
  wire [5:0] _sum_T_1 = $signed(man_buffer_two_complement_1) >>> exp_difference; // @[block_division.scala 287:15]
  wire [6:0] _sum_T_2 = $signed(man_buffer_two_complement_0) + $signed(_sum_T_1); // @[block_division.scala 285:46]
  wire [5:0] _sum_T_3 = $signed(man_buffer_two_complement_0) >>> exp_difference; // @[block_division.scala 290:15]
  wire [6:0] _sum_T_4 = $signed(man_buffer_two_complement_1) + $signed(_sum_T_3); // @[block_division.scala 288:50]
  wire [6:0] sum = _exp_buffer_0_T ? $signed(_sum_T_2) : $signed(_sum_T_4); // @[block_division.scala 283:24]
  wire [5:0] _man_buffer_two_complement_0_T_4 = ~sum[5:0]; // @[block_division.scala 292:78]
  wire [5:0] _man_buffer_two_complement_0_T_6 = _man_buffer_two_complement_0_T_4 + 6'h1; // @[block_division.scala 292:96]
  wire [5:0] _man_buffer_two_complement_0_T_8 = 6'h20 - 6'h1; // @[block_division.scala 292:116]
  wire [5:0] _man_buffer_two_complement_0_T_12 = 6'h1f - 6'h1; // @[block_division.scala 292:136]
  wire [5:0] _man_buffer_two_complement_0_T_14 = _man_buffer_two_complement_0_T_12 + 6'h1; // @[block_division.scala 292:143]
  wire [6:0] _man_buffer_two_complement_0_T_15 = _exp_buffer_0_T ? $signed(_sum_T_2) : $signed(_sum_T_4); // @[block_division.scala 292:154]
  wire [6:0] _man_buffer_two_complement_0_T_16 = _man_buffer_two_complement_0_T_6 > _man_buffer_two_complement_0_T_8 ?
    {{1'd0}, _man_buffer_two_complement_0_T_14} : _man_buffer_two_complement_0_T_15; // @[block_division.scala 292:75]
  wire [6:0] _man_buffer_two_complement_0_T_24 = sum[5:0] > _man_buffer_two_complement_0_T_8 ? {{1'd0},
    _man_buffer_two_complement_0_T_8} : _man_buffer_two_complement_0_T_15; // @[block_division.scala 293:14]
  wire [6:0] _man_buffer_two_complement_0_T_26 = sum[6] ? _man_buffer_two_complement_0_T_16 :
    _man_buffer_two_complement_0_T_24; // @[block_division.scala 293:83]
  wire  _exp_buffer_1_T = exp_buffer_2 > exp_buffer_3; // @[block_division.scala 274:31]
  wire [8:0] _exp_difference_T_7 = exp_buffer_2 - exp_buffer_3; // @[block_division.scala 280:31]
  wire [8:0] _exp_difference_T_9 = exp_buffer_3 - exp_buffer_2; // @[block_division.scala 281:35]
  wire [8:0] exp_difference_1 = _exp_buffer_1_T ? _exp_difference_T_7 : _exp_difference_T_9; // @[block_division.scala 278:35]
  wire [5:0] _sum_T_6 = $signed(man_buffer_two_complement_3) >>> exp_difference_1; // @[block_division.scala 287:15]
  wire [6:0] _sum_T_7 = $signed(man_buffer_two_complement_2) + $signed(_sum_T_6); // @[block_division.scala 285:46]
  wire [5:0] _sum_T_8 = $signed(man_buffer_two_complement_2) >>> exp_difference_1; // @[block_division.scala 290:15]
  wire [6:0] _sum_T_9 = $signed(man_buffer_two_complement_3) + $signed(_sum_T_8); // @[block_division.scala 288:50]
  wire [6:0] sum_1 = _exp_buffer_1_T ? $signed(_sum_T_7) : $signed(_sum_T_9); // @[block_division.scala 283:24]
  wire [5:0] _man_buffer_two_complement_1_T_4 = ~sum_1[5:0]; // @[block_division.scala 292:78]
  wire [5:0] _man_buffer_two_complement_1_T_6 = _man_buffer_two_complement_1_T_4 + 6'h1; // @[block_division.scala 292:96]
  wire [6:0] _man_buffer_two_complement_1_T_15 = _exp_buffer_1_T ? $signed(_sum_T_7) : $signed(_sum_T_9); // @[block_division.scala 292:154]
  wire [6:0] _man_buffer_two_complement_1_T_16 = _man_buffer_two_complement_1_T_6 > _man_buffer_two_complement_0_T_8 ?
    {{1'd0}, _man_buffer_two_complement_0_T_14} : _man_buffer_two_complement_1_T_15; // @[block_division.scala 292:75]
  wire [6:0] _man_buffer_two_complement_1_T_24 = sum_1[5:0] > _man_buffer_two_complement_0_T_8 ? {{1'd0},
    _man_buffer_two_complement_0_T_8} : _man_buffer_two_complement_1_T_15; // @[block_division.scala 293:14]
  wire [6:0] _man_buffer_two_complement_1_T_26 = sum_1[6] ? _man_buffer_two_complement_1_T_16 :
    _man_buffer_two_complement_1_T_24; // @[block_division.scala 293:83]
  wire [6:0] _GEN_13 = io_control_signal & enable ? $signed(_man_buffer_two_complement_0_T_26) : $signed({{1{_GEN_1[5
    ]}},_GEN_1}); // @[block_division.scala 266:47 292:40]
  wire [6:0] _GEN_15 = io_control_signal & enable ? $signed(_man_buffer_two_complement_1_T_26) : $signed({{1{_GEN_3[5
    ]}},_GEN_3}); // @[block_division.scala 266:47 292:40]
  reg [5:0] sign_man_hbfp; // @[block_division.scala 306:30]
  wire [5:0] _sign_man_hbfp_T_3 = {1'h0,man_buffer_two_complement_0[4:0]}; // @[block_division.scala 311:11]
  wire [5:0] _sign_man_hbfp_T_4 = ~_sign_man_hbfp_T_3; // @[block_division.scala 311:5]
  wire [5:0] _sign_man_hbfp_T_6 = _sign_man_hbfp_T_4 + 6'h1; // @[block_division.scala 311:60]
  wire [8:0] _io_result_tree_T_2 = {sign_man_hbfp[5],exp_buffer_0[8:1]}; // @[block_division.scala 329:38]
  wire [6:0] _GEN_17 = reset ? $signed(7'sh0) : $signed(_GEN_13); // @[block_division.scala 245:{12,12}]
  wire [6:0] _GEN_19 = reset ? $signed(7'sh0) : $signed(_GEN_15); // @[block_division.scala 245:{12,12}]
  assign io_result_tree = {_io_result_tree_T_2,sign_man_hbfp[4:0]}; // @[block_division.scala 329:61]
  always @(posedge clock) begin
    if (reset) begin // @[block_division.scala 243:60]
      exp_buffer_0 <= 9'h0; // @[block_division.scala 243:60]
    end else if (io_control_signal & enable) begin // @[block_division.scala 266:47]
      if (!(_exp_buffer_0_T)) begin // @[block_division.scala 273:33]
        exp_buffer_0 <= exp_buffer_1;
      end
    end else if (~io_control_signal) begin // @[block_division.scala 249:34]
      exp_buffer_0 <= io_exps_0; // @[block_division.scala 252:21]
    end
    if (reset) begin // @[block_division.scala 243:60]
      exp_buffer_1 <= 9'h0; // @[block_division.scala 243:60]
    end else if (io_control_signal & enable) begin // @[block_division.scala 266:47]
      if (_exp_buffer_1_T) begin // @[block_division.scala 273:33]
        exp_buffer_1 <= exp_buffer_2;
      end else begin
        exp_buffer_1 <= exp_buffer_3;
      end
    end else if (~io_control_signal) begin // @[block_division.scala 249:34]
      exp_buffer_1 <= io_exps_1; // @[block_division.scala 252:21]
    end
    if (reset) begin // @[block_division.scala 243:60]
      exp_buffer_2 <= 9'h0; // @[block_division.scala 243:60]
    end else if (~io_control_signal) begin // @[block_division.scala 249:34]
      exp_buffer_2 <= io_exps_2; // @[block_division.scala 252:21]
    end
    if (reset) begin // @[block_division.scala 243:60]
      exp_buffer_3 <= 9'h0; // @[block_division.scala 243:60]
    end else if (~io_control_signal) begin // @[block_division.scala 249:34]
      exp_buffer_3 <= io_exps_3; // @[block_division.scala 252:21]
    end
    man_buffer_two_complement_0 <= _GEN_17[5:0]; // @[block_division.scala 245:{12,12}]
    man_buffer_two_complement_1 <= _GEN_19[5:0]; // @[block_division.scala 245:{12,12}]
    if (reset) begin // @[block_division.scala 245:12]
      man_buffer_two_complement_2 <= 6'sh0; // @[block_division.scala 245:12]
    end else if (~io_control_signal) begin // @[block_division.scala 249:34]
      man_buffer_two_complement_2 <= io_sign_man_2; // @[block_division.scala 253:36]
    end
    if (reset) begin // @[block_division.scala 245:12]
      man_buffer_two_complement_3 <= 6'sh0; // @[block_division.scala 245:12]
    end else if (~io_control_signal) begin // @[block_division.scala 249:34]
      man_buffer_two_complement_3 <= io_sign_man_3; // @[block_division.scala 253:36]
    end
    if (reset) begin // @[block_division.scala 259:18]
      v <= 10'h0; // @[block_division.scala 259:18]
    end else if (io_control_signal & enable) begin // @[block_division.scala 266:47]
      v <= _v_T_1; // @[block_division.scala 270:11]
    end
    if (io_control_signal & enable) begin // @[block_division.scala 266:47]
      if (v == 10'h2) begin // @[block_division.scala 299:54]
        enable <= 1'h0; // @[block_division.scala 300:16]
      end else if (v == 10'h2) begin // @[block_division.scala 299:54]
        enable <= 1'h0; // @[block_division.scala 300:16]
      end else begin
        enable <= _GEN_8;
      end
    end else begin
      enable <= _GEN_8;
    end
    if (reset) begin // @[block_division.scala 306:30]
      sign_man_hbfp <= 6'h0; // @[block_division.scala 306:30]
    end else if (man_buffer_two_complement_0[5]) begin // @[block_division.scala 309:23]
      sign_man_hbfp <= _sign_man_hbfp_T_6;
    end else begin
      sign_man_hbfp <= man_buffer_two_complement_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  exp_buffer_0 = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  exp_buffer_1 = _RAND_1[8:0];
  _RAND_2 = {1{`RANDOM}};
  exp_buffer_2 = _RAND_2[8:0];
  _RAND_3 = {1{`RANDOM}};
  exp_buffer_3 = _RAND_3[8:0];
  _RAND_4 = {1{`RANDOM}};
  man_buffer_two_complement_0 = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  man_buffer_two_complement_1 = _RAND_5[5:0];
  _RAND_6 = {1{`RANDOM}};
  man_buffer_two_complement_2 = _RAND_6[5:0];
  _RAND_7 = {1{`RANDOM}};
  man_buffer_two_complement_3 = _RAND_7[5:0];
  _RAND_8 = {1{`RANDOM}};
  v = _RAND_8[9:0];
  _RAND_9 = {1{`RANDOM}};
  enable = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  sign_man_hbfp = _RAND_10[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module HbfpTensor(
  input         clock,
  input         reset,
  input  [4:0]  io_man_a_0,
  input  [4:0]  io_man_a_1,
  input  [4:0]  io_man_a_2,
  input  [4:0]  io_man_a_3,
  input  [4:0]  io_man_a_4,
  input  [4:0]  io_man_a_5,
  input  [4:0]  io_man_a_6,
  input  [4:0]  io_man_a_7,
  input  [4:0]  io_man_a_8,
  input  [4:0]  io_man_a_9,
  input  [4:0]  io_man_a_10,
  input  [4:0]  io_man_a_11,
  input  [4:0]  io_man_a_12,
  input  [4:0]  io_man_a_13,
  input  [4:0]  io_man_a_14,
  input  [4:0]  io_man_a_15,
  input  [4:0]  io_man_a_16,
  input  [4:0]  io_man_a_17,
  input  [4:0]  io_man_a_18,
  input  [4:0]  io_man_a_19,
  input  [4:0]  io_man_a_20,
  input  [4:0]  io_man_a_21,
  input  [4:0]  io_man_a_22,
  input  [4:0]  io_man_a_23,
  input  [4:0]  io_man_a_24,
  input  [4:0]  io_man_a_25,
  input  [4:0]  io_man_a_26,
  input  [4:0]  io_man_a_27,
  input  [4:0]  io_man_a_28,
  input  [4:0]  io_man_a_29,
  input  [4:0]  io_man_a_30,
  input  [4:0]  io_man_a_31,
  input  [4:0]  io_man_a_32,
  input  [4:0]  io_man_a_33,
  input  [4:0]  io_man_a_34,
  input  [4:0]  io_man_a_35,
  input  [4:0]  io_man_a_36,
  input  [4:0]  io_man_a_37,
  input  [4:0]  io_man_a_38,
  input  [4:0]  io_man_a_39,
  input  [4:0]  io_man_a_40,
  input  [4:0]  io_man_a_41,
  input  [4:0]  io_man_a_42,
  input  [4:0]  io_man_a_43,
  input  [4:0]  io_man_a_44,
  input  [4:0]  io_man_a_45,
  input  [4:0]  io_man_a_46,
  input  [4:0]  io_man_a_47,
  input  [4:0]  io_man_a_48,
  input  [4:0]  io_man_a_49,
  input  [4:0]  io_man_a_50,
  input  [4:0]  io_man_a_51,
  input  [4:0]  io_man_a_52,
  input  [4:0]  io_man_a_53,
  input  [4:0]  io_man_a_54,
  input  [4:0]  io_man_a_55,
  input  [4:0]  io_man_a_56,
  input  [4:0]  io_man_a_57,
  input  [4:0]  io_man_a_58,
  input  [4:0]  io_man_a_59,
  input  [4:0]  io_man_a_60,
  input  [4:0]  io_man_a_61,
  input  [4:0]  io_man_a_62,
  input  [4:0]  io_man_a_63,
  input  [4:0]  io_man_a_64,
  input  [4:0]  io_man_a_65,
  input  [4:0]  io_man_a_66,
  input  [4:0]  io_man_a_67,
  input  [4:0]  io_man_a_68,
  input  [4:0]  io_man_a_69,
  input  [4:0]  io_man_a_70,
  input  [4:0]  io_man_a_71,
  input  [4:0]  io_man_a_72,
  input  [4:0]  io_man_a_73,
  input  [4:0]  io_man_a_74,
  input  [4:0]  io_man_a_75,
  input  [4:0]  io_man_a_76,
  input  [4:0]  io_man_a_77,
  input  [4:0]  io_man_a_78,
  input  [4:0]  io_man_a_79,
  input  [4:0]  io_man_a_80,
  input  [4:0]  io_man_a_81,
  input  [4:0]  io_man_a_82,
  input  [4:0]  io_man_a_83,
  input  [4:0]  io_man_a_84,
  input  [4:0]  io_man_a_85,
  input  [4:0]  io_man_a_86,
  input  [4:0]  io_man_a_87,
  input  [4:0]  io_man_a_88,
  input  [4:0]  io_man_a_89,
  input  [4:0]  io_man_a_90,
  input  [4:0]  io_man_a_91,
  input  [4:0]  io_man_a_92,
  input  [4:0]  io_man_a_93,
  input  [4:0]  io_man_a_94,
  input  [4:0]  io_man_a_95,
  input  [4:0]  io_man_a_96,
  input  [4:0]  io_man_a_97,
  input  [4:0]  io_man_a_98,
  input  [4:0]  io_man_a_99,
  input  [4:0]  io_man_a_100,
  input  [4:0]  io_man_a_101,
  input  [4:0]  io_man_a_102,
  input  [4:0]  io_man_a_103,
  input  [4:0]  io_man_a_104,
  input  [4:0]  io_man_a_105,
  input  [4:0]  io_man_a_106,
  input  [4:0]  io_man_a_107,
  input  [4:0]  io_man_a_108,
  input  [4:0]  io_man_a_109,
  input  [4:0]  io_man_a_110,
  input  [4:0]  io_man_a_111,
  input  [4:0]  io_man_a_112,
  input  [4:0]  io_man_a_113,
  input  [4:0]  io_man_a_114,
  input  [4:0]  io_man_a_115,
  input  [4:0]  io_man_a_116,
  input  [4:0]  io_man_a_117,
  input  [4:0]  io_man_a_118,
  input  [4:0]  io_man_a_119,
  input  [4:0]  io_man_a_120,
  input  [4:0]  io_man_a_121,
  input  [4:0]  io_man_a_122,
  input  [4:0]  io_man_a_123,
  input  [4:0]  io_man_a_124,
  input  [4:0]  io_man_a_125,
  input  [4:0]  io_man_a_126,
  input  [4:0]  io_man_a_127,
  input  [4:0]  io_man_a_128,
  input  [4:0]  io_man_a_129,
  input  [4:0]  io_man_a_130,
  input  [4:0]  io_man_a_131,
  input  [4:0]  io_man_a_132,
  input  [4:0]  io_man_a_133,
  input  [4:0]  io_man_a_134,
  input  [4:0]  io_man_a_135,
  input  [4:0]  io_man_a_136,
  input  [4:0]  io_man_a_137,
  input  [4:0]  io_man_a_138,
  input  [4:0]  io_man_a_139,
  input  [4:0]  io_man_a_140,
  input  [4:0]  io_man_a_141,
  input  [4:0]  io_man_a_142,
  input  [4:0]  io_man_a_143,
  input  [4:0]  io_man_a_144,
  input  [4:0]  io_man_a_145,
  input  [4:0]  io_man_a_146,
  input  [4:0]  io_man_a_147,
  input  [4:0]  io_man_a_148,
  input  [4:0]  io_man_a_149,
  input  [4:0]  io_man_a_150,
  input  [4:0]  io_man_a_151,
  input  [4:0]  io_man_a_152,
  input  [4:0]  io_man_a_153,
  input  [4:0]  io_man_a_154,
  input  [4:0]  io_man_a_155,
  input  [4:0]  io_man_a_156,
  input  [4:0]  io_man_a_157,
  input  [4:0]  io_man_a_158,
  input  [4:0]  io_man_a_159,
  input  [4:0]  io_man_a_160,
  input  [4:0]  io_man_a_161,
  input  [4:0]  io_man_a_162,
  input  [4:0]  io_man_a_163,
  input  [4:0]  io_man_a_164,
  input  [4:0]  io_man_a_165,
  input  [4:0]  io_man_a_166,
  input  [4:0]  io_man_a_167,
  input  [4:0]  io_man_a_168,
  input  [4:0]  io_man_a_169,
  input  [4:0]  io_man_a_170,
  input  [4:0]  io_man_a_171,
  input  [4:0]  io_man_a_172,
  input  [4:0]  io_man_a_173,
  input  [4:0]  io_man_a_174,
  input  [4:0]  io_man_a_175,
  input  [4:0]  io_man_a_176,
  input  [4:0]  io_man_a_177,
  input  [4:0]  io_man_a_178,
  input  [4:0]  io_man_a_179,
  input  [4:0]  io_man_a_180,
  input  [4:0]  io_man_a_181,
  input  [4:0]  io_man_a_182,
  input  [4:0]  io_man_a_183,
  input  [4:0]  io_man_a_184,
  input  [4:0]  io_man_a_185,
  input  [4:0]  io_man_a_186,
  input  [4:0]  io_man_a_187,
  input  [4:0]  io_man_a_188,
  input  [4:0]  io_man_a_189,
  input  [4:0]  io_man_a_190,
  input  [4:0]  io_man_a_191,
  input  [4:0]  io_man_a_192,
  input  [4:0]  io_man_a_193,
  input  [4:0]  io_man_a_194,
  input  [4:0]  io_man_a_195,
  input  [4:0]  io_man_a_196,
  input  [4:0]  io_man_a_197,
  input  [4:0]  io_man_a_198,
  input  [4:0]  io_man_a_199,
  input  [4:0]  io_man_a_200,
  input  [4:0]  io_man_a_201,
  input  [4:0]  io_man_a_202,
  input  [4:0]  io_man_a_203,
  input  [4:0]  io_man_a_204,
  input  [4:0]  io_man_a_205,
  input  [4:0]  io_man_a_206,
  input  [4:0]  io_man_a_207,
  input  [4:0]  io_man_a_208,
  input  [4:0]  io_man_a_209,
  input  [4:0]  io_man_a_210,
  input  [4:0]  io_man_a_211,
  input  [4:0]  io_man_a_212,
  input  [4:0]  io_man_a_213,
  input  [4:0]  io_man_a_214,
  input  [4:0]  io_man_a_215,
  input  [4:0]  io_man_a_216,
  input  [4:0]  io_man_a_217,
  input  [4:0]  io_man_a_218,
  input  [4:0]  io_man_a_219,
  input  [4:0]  io_man_a_220,
  input  [4:0]  io_man_a_221,
  input  [4:0]  io_man_a_222,
  input  [4:0]  io_man_a_223,
  input  [4:0]  io_man_a_224,
  input  [4:0]  io_man_a_225,
  input  [4:0]  io_man_a_226,
  input  [4:0]  io_man_a_227,
  input  [4:0]  io_man_a_228,
  input  [4:0]  io_man_a_229,
  input  [4:0]  io_man_a_230,
  input  [4:0]  io_man_a_231,
  input  [4:0]  io_man_a_232,
  input  [4:0]  io_man_a_233,
  input  [4:0]  io_man_a_234,
  input  [4:0]  io_man_a_235,
  input  [4:0]  io_man_a_236,
  input  [4:0]  io_man_a_237,
  input  [4:0]  io_man_a_238,
  input  [4:0]  io_man_a_239,
  input  [4:0]  io_man_a_240,
  input  [4:0]  io_man_a_241,
  input  [4:0]  io_man_a_242,
  input  [4:0]  io_man_a_243,
  input  [4:0]  io_man_a_244,
  input  [4:0]  io_man_a_245,
  input  [4:0]  io_man_a_246,
  input  [4:0]  io_man_a_247,
  input  [4:0]  io_man_a_248,
  input  [4:0]  io_man_a_249,
  input  [4:0]  io_man_a_250,
  input  [4:0]  io_man_a_251,
  input  [4:0]  io_man_a_252,
  input  [4:0]  io_man_a_253,
  input  [4:0]  io_man_a_254,
  input  [4:0]  io_man_a_255,
  input  [4:0]  io_man_b_0,
  input  [4:0]  io_man_b_1,
  input  [4:0]  io_man_b_2,
  input  [4:0]  io_man_b_3,
  input  [4:0]  io_man_b_4,
  input  [4:0]  io_man_b_5,
  input  [4:0]  io_man_b_6,
  input  [4:0]  io_man_b_7,
  input  [4:0]  io_man_b_8,
  input  [4:0]  io_man_b_9,
  input  [4:0]  io_man_b_10,
  input  [4:0]  io_man_b_11,
  input  [4:0]  io_man_b_12,
  input  [4:0]  io_man_b_13,
  input  [4:0]  io_man_b_14,
  input  [4:0]  io_man_b_15,
  input  [4:0]  io_man_b_16,
  input  [4:0]  io_man_b_17,
  input  [4:0]  io_man_b_18,
  input  [4:0]  io_man_b_19,
  input  [4:0]  io_man_b_20,
  input  [4:0]  io_man_b_21,
  input  [4:0]  io_man_b_22,
  input  [4:0]  io_man_b_23,
  input  [4:0]  io_man_b_24,
  input  [4:0]  io_man_b_25,
  input  [4:0]  io_man_b_26,
  input  [4:0]  io_man_b_27,
  input  [4:0]  io_man_b_28,
  input  [4:0]  io_man_b_29,
  input  [4:0]  io_man_b_30,
  input  [4:0]  io_man_b_31,
  input  [4:0]  io_man_b_32,
  input  [4:0]  io_man_b_33,
  input  [4:0]  io_man_b_34,
  input  [4:0]  io_man_b_35,
  input  [4:0]  io_man_b_36,
  input  [4:0]  io_man_b_37,
  input  [4:0]  io_man_b_38,
  input  [4:0]  io_man_b_39,
  input  [4:0]  io_man_b_40,
  input  [4:0]  io_man_b_41,
  input  [4:0]  io_man_b_42,
  input  [4:0]  io_man_b_43,
  input  [4:0]  io_man_b_44,
  input  [4:0]  io_man_b_45,
  input  [4:0]  io_man_b_46,
  input  [4:0]  io_man_b_47,
  input  [4:0]  io_man_b_48,
  input  [4:0]  io_man_b_49,
  input  [4:0]  io_man_b_50,
  input  [4:0]  io_man_b_51,
  input  [4:0]  io_man_b_52,
  input  [4:0]  io_man_b_53,
  input  [4:0]  io_man_b_54,
  input  [4:0]  io_man_b_55,
  input  [4:0]  io_man_b_56,
  input  [4:0]  io_man_b_57,
  input  [4:0]  io_man_b_58,
  input  [4:0]  io_man_b_59,
  input  [4:0]  io_man_b_60,
  input  [4:0]  io_man_b_61,
  input  [4:0]  io_man_b_62,
  input  [4:0]  io_man_b_63,
  input  [4:0]  io_man_b_64,
  input  [4:0]  io_man_b_65,
  input  [4:0]  io_man_b_66,
  input  [4:0]  io_man_b_67,
  input  [4:0]  io_man_b_68,
  input  [4:0]  io_man_b_69,
  input  [4:0]  io_man_b_70,
  input  [4:0]  io_man_b_71,
  input  [4:0]  io_man_b_72,
  input  [4:0]  io_man_b_73,
  input  [4:0]  io_man_b_74,
  input  [4:0]  io_man_b_75,
  input  [4:0]  io_man_b_76,
  input  [4:0]  io_man_b_77,
  input  [4:0]  io_man_b_78,
  input  [4:0]  io_man_b_79,
  input  [4:0]  io_man_b_80,
  input  [4:0]  io_man_b_81,
  input  [4:0]  io_man_b_82,
  input  [4:0]  io_man_b_83,
  input  [4:0]  io_man_b_84,
  input  [4:0]  io_man_b_85,
  input  [4:0]  io_man_b_86,
  input  [4:0]  io_man_b_87,
  input  [4:0]  io_man_b_88,
  input  [4:0]  io_man_b_89,
  input  [4:0]  io_man_b_90,
  input  [4:0]  io_man_b_91,
  input  [4:0]  io_man_b_92,
  input  [4:0]  io_man_b_93,
  input  [4:0]  io_man_b_94,
  input  [4:0]  io_man_b_95,
  input  [4:0]  io_man_b_96,
  input  [4:0]  io_man_b_97,
  input  [4:0]  io_man_b_98,
  input  [4:0]  io_man_b_99,
  input  [4:0]  io_man_b_100,
  input  [4:0]  io_man_b_101,
  input  [4:0]  io_man_b_102,
  input  [4:0]  io_man_b_103,
  input  [4:0]  io_man_b_104,
  input  [4:0]  io_man_b_105,
  input  [4:0]  io_man_b_106,
  input  [4:0]  io_man_b_107,
  input  [4:0]  io_man_b_108,
  input  [4:0]  io_man_b_109,
  input  [4:0]  io_man_b_110,
  input  [4:0]  io_man_b_111,
  input  [4:0]  io_man_b_112,
  input  [4:0]  io_man_b_113,
  input  [4:0]  io_man_b_114,
  input  [4:0]  io_man_b_115,
  input  [4:0]  io_man_b_116,
  input  [4:0]  io_man_b_117,
  input  [4:0]  io_man_b_118,
  input  [4:0]  io_man_b_119,
  input  [4:0]  io_man_b_120,
  input  [4:0]  io_man_b_121,
  input  [4:0]  io_man_b_122,
  input  [4:0]  io_man_b_123,
  input  [4:0]  io_man_b_124,
  input  [4:0]  io_man_b_125,
  input  [4:0]  io_man_b_126,
  input  [4:0]  io_man_b_127,
  input  [4:0]  io_man_b_128,
  input  [4:0]  io_man_b_129,
  input  [4:0]  io_man_b_130,
  input  [4:0]  io_man_b_131,
  input  [4:0]  io_man_b_132,
  input  [4:0]  io_man_b_133,
  input  [4:0]  io_man_b_134,
  input  [4:0]  io_man_b_135,
  input  [4:0]  io_man_b_136,
  input  [4:0]  io_man_b_137,
  input  [4:0]  io_man_b_138,
  input  [4:0]  io_man_b_139,
  input  [4:0]  io_man_b_140,
  input  [4:0]  io_man_b_141,
  input  [4:0]  io_man_b_142,
  input  [4:0]  io_man_b_143,
  input  [4:0]  io_man_b_144,
  input  [4:0]  io_man_b_145,
  input  [4:0]  io_man_b_146,
  input  [4:0]  io_man_b_147,
  input  [4:0]  io_man_b_148,
  input  [4:0]  io_man_b_149,
  input  [4:0]  io_man_b_150,
  input  [4:0]  io_man_b_151,
  input  [4:0]  io_man_b_152,
  input  [4:0]  io_man_b_153,
  input  [4:0]  io_man_b_154,
  input  [4:0]  io_man_b_155,
  input  [4:0]  io_man_b_156,
  input  [4:0]  io_man_b_157,
  input  [4:0]  io_man_b_158,
  input  [4:0]  io_man_b_159,
  input  [4:0]  io_man_b_160,
  input  [4:0]  io_man_b_161,
  input  [4:0]  io_man_b_162,
  input  [4:0]  io_man_b_163,
  input  [4:0]  io_man_b_164,
  input  [4:0]  io_man_b_165,
  input  [4:0]  io_man_b_166,
  input  [4:0]  io_man_b_167,
  input  [4:0]  io_man_b_168,
  input  [4:0]  io_man_b_169,
  input  [4:0]  io_man_b_170,
  input  [4:0]  io_man_b_171,
  input  [4:0]  io_man_b_172,
  input  [4:0]  io_man_b_173,
  input  [4:0]  io_man_b_174,
  input  [4:0]  io_man_b_175,
  input  [4:0]  io_man_b_176,
  input  [4:0]  io_man_b_177,
  input  [4:0]  io_man_b_178,
  input  [4:0]  io_man_b_179,
  input  [4:0]  io_man_b_180,
  input  [4:0]  io_man_b_181,
  input  [4:0]  io_man_b_182,
  input  [4:0]  io_man_b_183,
  input  [4:0]  io_man_b_184,
  input  [4:0]  io_man_b_185,
  input  [4:0]  io_man_b_186,
  input  [4:0]  io_man_b_187,
  input  [4:0]  io_man_b_188,
  input  [4:0]  io_man_b_189,
  input  [4:0]  io_man_b_190,
  input  [4:0]  io_man_b_191,
  input  [4:0]  io_man_b_192,
  input  [4:0]  io_man_b_193,
  input  [4:0]  io_man_b_194,
  input  [4:0]  io_man_b_195,
  input  [4:0]  io_man_b_196,
  input  [4:0]  io_man_b_197,
  input  [4:0]  io_man_b_198,
  input  [4:0]  io_man_b_199,
  input  [4:0]  io_man_b_200,
  input  [4:0]  io_man_b_201,
  input  [4:0]  io_man_b_202,
  input  [4:0]  io_man_b_203,
  input  [4:0]  io_man_b_204,
  input  [4:0]  io_man_b_205,
  input  [4:0]  io_man_b_206,
  input  [4:0]  io_man_b_207,
  input  [4:0]  io_man_b_208,
  input  [4:0]  io_man_b_209,
  input  [4:0]  io_man_b_210,
  input  [4:0]  io_man_b_211,
  input  [4:0]  io_man_b_212,
  input  [4:0]  io_man_b_213,
  input  [4:0]  io_man_b_214,
  input  [4:0]  io_man_b_215,
  input  [4:0]  io_man_b_216,
  input  [4:0]  io_man_b_217,
  input  [4:0]  io_man_b_218,
  input  [4:0]  io_man_b_219,
  input  [4:0]  io_man_b_220,
  input  [4:0]  io_man_b_221,
  input  [4:0]  io_man_b_222,
  input  [4:0]  io_man_b_223,
  input  [4:0]  io_man_b_224,
  input  [4:0]  io_man_b_225,
  input  [4:0]  io_man_b_226,
  input  [4:0]  io_man_b_227,
  input  [4:0]  io_man_b_228,
  input  [4:0]  io_man_b_229,
  input  [4:0]  io_man_b_230,
  input  [4:0]  io_man_b_231,
  input  [4:0]  io_man_b_232,
  input  [4:0]  io_man_b_233,
  input  [4:0]  io_man_b_234,
  input  [4:0]  io_man_b_235,
  input  [4:0]  io_man_b_236,
  input  [4:0]  io_man_b_237,
  input  [4:0]  io_man_b_238,
  input  [4:0]  io_man_b_239,
  input  [4:0]  io_man_b_240,
  input  [4:0]  io_man_b_241,
  input  [4:0]  io_man_b_242,
  input  [4:0]  io_man_b_243,
  input  [4:0]  io_man_b_244,
  input  [4:0]  io_man_b_245,
  input  [4:0]  io_man_b_246,
  input  [4:0]  io_man_b_247,
  input  [4:0]  io_man_b_248,
  input  [4:0]  io_man_b_249,
  input  [4:0]  io_man_b_250,
  input  [4:0]  io_man_b_251,
  input  [4:0]  io_man_b_252,
  input  [4:0]  io_man_b_253,
  input  [4:0]  io_man_b_254,
  input  [4:0]  io_man_b_255,
  input         io_sign_a_0,
  input         io_sign_a_1,
  input         io_sign_a_2,
  input         io_sign_a_3,
  input         io_sign_a_4,
  input         io_sign_a_5,
  input         io_sign_a_6,
  input         io_sign_a_7,
  input         io_sign_a_8,
  input         io_sign_a_9,
  input         io_sign_a_10,
  input         io_sign_a_11,
  input         io_sign_a_12,
  input         io_sign_a_13,
  input         io_sign_a_14,
  input         io_sign_a_15,
  input         io_sign_a_16,
  input         io_sign_a_17,
  input         io_sign_a_18,
  input         io_sign_a_19,
  input         io_sign_a_20,
  input         io_sign_a_21,
  input         io_sign_a_22,
  input         io_sign_a_23,
  input         io_sign_a_24,
  input         io_sign_a_25,
  input         io_sign_a_26,
  input         io_sign_a_27,
  input         io_sign_a_28,
  input         io_sign_a_29,
  input         io_sign_a_30,
  input         io_sign_a_31,
  input         io_sign_a_32,
  input         io_sign_a_33,
  input         io_sign_a_34,
  input         io_sign_a_35,
  input         io_sign_a_36,
  input         io_sign_a_37,
  input         io_sign_a_38,
  input         io_sign_a_39,
  input         io_sign_a_40,
  input         io_sign_a_41,
  input         io_sign_a_42,
  input         io_sign_a_43,
  input         io_sign_a_44,
  input         io_sign_a_45,
  input         io_sign_a_46,
  input         io_sign_a_47,
  input         io_sign_a_48,
  input         io_sign_a_49,
  input         io_sign_a_50,
  input         io_sign_a_51,
  input         io_sign_a_52,
  input         io_sign_a_53,
  input         io_sign_a_54,
  input         io_sign_a_55,
  input         io_sign_a_56,
  input         io_sign_a_57,
  input         io_sign_a_58,
  input         io_sign_a_59,
  input         io_sign_a_60,
  input         io_sign_a_61,
  input         io_sign_a_62,
  input         io_sign_a_63,
  input         io_sign_a_64,
  input         io_sign_a_65,
  input         io_sign_a_66,
  input         io_sign_a_67,
  input         io_sign_a_68,
  input         io_sign_a_69,
  input         io_sign_a_70,
  input         io_sign_a_71,
  input         io_sign_a_72,
  input         io_sign_a_73,
  input         io_sign_a_74,
  input         io_sign_a_75,
  input         io_sign_a_76,
  input         io_sign_a_77,
  input         io_sign_a_78,
  input         io_sign_a_79,
  input         io_sign_a_80,
  input         io_sign_a_81,
  input         io_sign_a_82,
  input         io_sign_a_83,
  input         io_sign_a_84,
  input         io_sign_a_85,
  input         io_sign_a_86,
  input         io_sign_a_87,
  input         io_sign_a_88,
  input         io_sign_a_89,
  input         io_sign_a_90,
  input         io_sign_a_91,
  input         io_sign_a_92,
  input         io_sign_a_93,
  input         io_sign_a_94,
  input         io_sign_a_95,
  input         io_sign_a_96,
  input         io_sign_a_97,
  input         io_sign_a_98,
  input         io_sign_a_99,
  input         io_sign_a_100,
  input         io_sign_a_101,
  input         io_sign_a_102,
  input         io_sign_a_103,
  input         io_sign_a_104,
  input         io_sign_a_105,
  input         io_sign_a_106,
  input         io_sign_a_107,
  input         io_sign_a_108,
  input         io_sign_a_109,
  input         io_sign_a_110,
  input         io_sign_a_111,
  input         io_sign_a_112,
  input         io_sign_a_113,
  input         io_sign_a_114,
  input         io_sign_a_115,
  input         io_sign_a_116,
  input         io_sign_a_117,
  input         io_sign_a_118,
  input         io_sign_a_119,
  input         io_sign_a_120,
  input         io_sign_a_121,
  input         io_sign_a_122,
  input         io_sign_a_123,
  input         io_sign_a_124,
  input         io_sign_a_125,
  input         io_sign_a_126,
  input         io_sign_a_127,
  input         io_sign_a_128,
  input         io_sign_a_129,
  input         io_sign_a_130,
  input         io_sign_a_131,
  input         io_sign_a_132,
  input         io_sign_a_133,
  input         io_sign_a_134,
  input         io_sign_a_135,
  input         io_sign_a_136,
  input         io_sign_a_137,
  input         io_sign_a_138,
  input         io_sign_a_139,
  input         io_sign_a_140,
  input         io_sign_a_141,
  input         io_sign_a_142,
  input         io_sign_a_143,
  input         io_sign_a_144,
  input         io_sign_a_145,
  input         io_sign_a_146,
  input         io_sign_a_147,
  input         io_sign_a_148,
  input         io_sign_a_149,
  input         io_sign_a_150,
  input         io_sign_a_151,
  input         io_sign_a_152,
  input         io_sign_a_153,
  input         io_sign_a_154,
  input         io_sign_a_155,
  input         io_sign_a_156,
  input         io_sign_a_157,
  input         io_sign_a_158,
  input         io_sign_a_159,
  input         io_sign_a_160,
  input         io_sign_a_161,
  input         io_sign_a_162,
  input         io_sign_a_163,
  input         io_sign_a_164,
  input         io_sign_a_165,
  input         io_sign_a_166,
  input         io_sign_a_167,
  input         io_sign_a_168,
  input         io_sign_a_169,
  input         io_sign_a_170,
  input         io_sign_a_171,
  input         io_sign_a_172,
  input         io_sign_a_173,
  input         io_sign_a_174,
  input         io_sign_a_175,
  input         io_sign_a_176,
  input         io_sign_a_177,
  input         io_sign_a_178,
  input         io_sign_a_179,
  input         io_sign_a_180,
  input         io_sign_a_181,
  input         io_sign_a_182,
  input         io_sign_a_183,
  input         io_sign_a_184,
  input         io_sign_a_185,
  input         io_sign_a_186,
  input         io_sign_a_187,
  input         io_sign_a_188,
  input         io_sign_a_189,
  input         io_sign_a_190,
  input         io_sign_a_191,
  input         io_sign_a_192,
  input         io_sign_a_193,
  input         io_sign_a_194,
  input         io_sign_a_195,
  input         io_sign_a_196,
  input         io_sign_a_197,
  input         io_sign_a_198,
  input         io_sign_a_199,
  input         io_sign_a_200,
  input         io_sign_a_201,
  input         io_sign_a_202,
  input         io_sign_a_203,
  input         io_sign_a_204,
  input         io_sign_a_205,
  input         io_sign_a_206,
  input         io_sign_a_207,
  input         io_sign_a_208,
  input         io_sign_a_209,
  input         io_sign_a_210,
  input         io_sign_a_211,
  input         io_sign_a_212,
  input         io_sign_a_213,
  input         io_sign_a_214,
  input         io_sign_a_215,
  input         io_sign_a_216,
  input         io_sign_a_217,
  input         io_sign_a_218,
  input         io_sign_a_219,
  input         io_sign_a_220,
  input         io_sign_a_221,
  input         io_sign_a_222,
  input         io_sign_a_223,
  input         io_sign_a_224,
  input         io_sign_a_225,
  input         io_sign_a_226,
  input         io_sign_a_227,
  input         io_sign_a_228,
  input         io_sign_a_229,
  input         io_sign_a_230,
  input         io_sign_a_231,
  input         io_sign_a_232,
  input         io_sign_a_233,
  input         io_sign_a_234,
  input         io_sign_a_235,
  input         io_sign_a_236,
  input         io_sign_a_237,
  input         io_sign_a_238,
  input         io_sign_a_239,
  input         io_sign_a_240,
  input         io_sign_a_241,
  input         io_sign_a_242,
  input         io_sign_a_243,
  input         io_sign_a_244,
  input         io_sign_a_245,
  input         io_sign_a_246,
  input         io_sign_a_247,
  input         io_sign_a_248,
  input         io_sign_a_249,
  input         io_sign_a_250,
  input         io_sign_a_251,
  input         io_sign_a_252,
  input         io_sign_a_253,
  input         io_sign_a_254,
  input         io_sign_a_255,
  input         io_sign_b_0,
  input         io_sign_b_1,
  input         io_sign_b_2,
  input         io_sign_b_3,
  input         io_sign_b_4,
  input         io_sign_b_5,
  input         io_sign_b_6,
  input         io_sign_b_7,
  input         io_sign_b_8,
  input         io_sign_b_9,
  input         io_sign_b_10,
  input         io_sign_b_11,
  input         io_sign_b_12,
  input         io_sign_b_13,
  input         io_sign_b_14,
  input         io_sign_b_15,
  input         io_sign_b_16,
  input         io_sign_b_17,
  input         io_sign_b_18,
  input         io_sign_b_19,
  input         io_sign_b_20,
  input         io_sign_b_21,
  input         io_sign_b_22,
  input         io_sign_b_23,
  input         io_sign_b_24,
  input         io_sign_b_25,
  input         io_sign_b_26,
  input         io_sign_b_27,
  input         io_sign_b_28,
  input         io_sign_b_29,
  input         io_sign_b_30,
  input         io_sign_b_31,
  input         io_sign_b_32,
  input         io_sign_b_33,
  input         io_sign_b_34,
  input         io_sign_b_35,
  input         io_sign_b_36,
  input         io_sign_b_37,
  input         io_sign_b_38,
  input         io_sign_b_39,
  input         io_sign_b_40,
  input         io_sign_b_41,
  input         io_sign_b_42,
  input         io_sign_b_43,
  input         io_sign_b_44,
  input         io_sign_b_45,
  input         io_sign_b_46,
  input         io_sign_b_47,
  input         io_sign_b_48,
  input         io_sign_b_49,
  input         io_sign_b_50,
  input         io_sign_b_51,
  input         io_sign_b_52,
  input         io_sign_b_53,
  input         io_sign_b_54,
  input         io_sign_b_55,
  input         io_sign_b_56,
  input         io_sign_b_57,
  input         io_sign_b_58,
  input         io_sign_b_59,
  input         io_sign_b_60,
  input         io_sign_b_61,
  input         io_sign_b_62,
  input         io_sign_b_63,
  input         io_sign_b_64,
  input         io_sign_b_65,
  input         io_sign_b_66,
  input         io_sign_b_67,
  input         io_sign_b_68,
  input         io_sign_b_69,
  input         io_sign_b_70,
  input         io_sign_b_71,
  input         io_sign_b_72,
  input         io_sign_b_73,
  input         io_sign_b_74,
  input         io_sign_b_75,
  input         io_sign_b_76,
  input         io_sign_b_77,
  input         io_sign_b_78,
  input         io_sign_b_79,
  input         io_sign_b_80,
  input         io_sign_b_81,
  input         io_sign_b_82,
  input         io_sign_b_83,
  input         io_sign_b_84,
  input         io_sign_b_85,
  input         io_sign_b_86,
  input         io_sign_b_87,
  input         io_sign_b_88,
  input         io_sign_b_89,
  input         io_sign_b_90,
  input         io_sign_b_91,
  input         io_sign_b_92,
  input         io_sign_b_93,
  input         io_sign_b_94,
  input         io_sign_b_95,
  input         io_sign_b_96,
  input         io_sign_b_97,
  input         io_sign_b_98,
  input         io_sign_b_99,
  input         io_sign_b_100,
  input         io_sign_b_101,
  input         io_sign_b_102,
  input         io_sign_b_103,
  input         io_sign_b_104,
  input         io_sign_b_105,
  input         io_sign_b_106,
  input         io_sign_b_107,
  input         io_sign_b_108,
  input         io_sign_b_109,
  input         io_sign_b_110,
  input         io_sign_b_111,
  input         io_sign_b_112,
  input         io_sign_b_113,
  input         io_sign_b_114,
  input         io_sign_b_115,
  input         io_sign_b_116,
  input         io_sign_b_117,
  input         io_sign_b_118,
  input         io_sign_b_119,
  input         io_sign_b_120,
  input         io_sign_b_121,
  input         io_sign_b_122,
  input         io_sign_b_123,
  input         io_sign_b_124,
  input         io_sign_b_125,
  input         io_sign_b_126,
  input         io_sign_b_127,
  input         io_sign_b_128,
  input         io_sign_b_129,
  input         io_sign_b_130,
  input         io_sign_b_131,
  input         io_sign_b_132,
  input         io_sign_b_133,
  input         io_sign_b_134,
  input         io_sign_b_135,
  input         io_sign_b_136,
  input         io_sign_b_137,
  input         io_sign_b_138,
  input         io_sign_b_139,
  input         io_sign_b_140,
  input         io_sign_b_141,
  input         io_sign_b_142,
  input         io_sign_b_143,
  input         io_sign_b_144,
  input         io_sign_b_145,
  input         io_sign_b_146,
  input         io_sign_b_147,
  input         io_sign_b_148,
  input         io_sign_b_149,
  input         io_sign_b_150,
  input         io_sign_b_151,
  input         io_sign_b_152,
  input         io_sign_b_153,
  input         io_sign_b_154,
  input         io_sign_b_155,
  input         io_sign_b_156,
  input         io_sign_b_157,
  input         io_sign_b_158,
  input         io_sign_b_159,
  input         io_sign_b_160,
  input         io_sign_b_161,
  input         io_sign_b_162,
  input         io_sign_b_163,
  input         io_sign_b_164,
  input         io_sign_b_165,
  input         io_sign_b_166,
  input         io_sign_b_167,
  input         io_sign_b_168,
  input         io_sign_b_169,
  input         io_sign_b_170,
  input         io_sign_b_171,
  input         io_sign_b_172,
  input         io_sign_b_173,
  input         io_sign_b_174,
  input         io_sign_b_175,
  input         io_sign_b_176,
  input         io_sign_b_177,
  input         io_sign_b_178,
  input         io_sign_b_179,
  input         io_sign_b_180,
  input         io_sign_b_181,
  input         io_sign_b_182,
  input         io_sign_b_183,
  input         io_sign_b_184,
  input         io_sign_b_185,
  input         io_sign_b_186,
  input         io_sign_b_187,
  input         io_sign_b_188,
  input         io_sign_b_189,
  input         io_sign_b_190,
  input         io_sign_b_191,
  input         io_sign_b_192,
  input         io_sign_b_193,
  input         io_sign_b_194,
  input         io_sign_b_195,
  input         io_sign_b_196,
  input         io_sign_b_197,
  input         io_sign_b_198,
  input         io_sign_b_199,
  input         io_sign_b_200,
  input         io_sign_b_201,
  input         io_sign_b_202,
  input         io_sign_b_203,
  input         io_sign_b_204,
  input         io_sign_b_205,
  input         io_sign_b_206,
  input         io_sign_b_207,
  input         io_sign_b_208,
  input         io_sign_b_209,
  input         io_sign_b_210,
  input         io_sign_b_211,
  input         io_sign_b_212,
  input         io_sign_b_213,
  input         io_sign_b_214,
  input         io_sign_b_215,
  input         io_sign_b_216,
  input         io_sign_b_217,
  input         io_sign_b_218,
  input         io_sign_b_219,
  input         io_sign_b_220,
  input         io_sign_b_221,
  input         io_sign_b_222,
  input         io_sign_b_223,
  input         io_sign_b_224,
  input         io_sign_b_225,
  input         io_sign_b_226,
  input         io_sign_b_227,
  input         io_sign_b_228,
  input         io_sign_b_229,
  input         io_sign_b_230,
  input         io_sign_b_231,
  input         io_sign_b_232,
  input         io_sign_b_233,
  input         io_sign_b_234,
  input         io_sign_b_235,
  input         io_sign_b_236,
  input         io_sign_b_237,
  input         io_sign_b_238,
  input         io_sign_b_239,
  input         io_sign_b_240,
  input         io_sign_b_241,
  input         io_sign_b_242,
  input         io_sign_b_243,
  input         io_sign_b_244,
  input         io_sign_b_245,
  input         io_sign_b_246,
  input         io_sign_b_247,
  input         io_sign_b_248,
  input         io_sign_b_249,
  input         io_sign_b_250,
  input         io_sign_b_251,
  input         io_sign_b_252,
  input         io_sign_b_253,
  input         io_sign_b_254,
  input         io_sign_b_255,
  input  [7:0]  io_exp_a_0,
  input  [7:0]  io_exp_a_1,
  input  [7:0]  io_exp_a_2,
  input  [7:0]  io_exp_a_3,
  input  [7:0]  io_exp_b_0,
  input  [7:0]  io_exp_b_1,
  input  [7:0]  io_exp_b_2,
  input  [7:0]  io_exp_b_3,
  input         io_control,
  input         io_control2,
  output [13:0] io_result
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1305;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1329;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [31:0] _RAND_1334;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [31:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1377;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [31:0] _RAND_1413;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1434;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1461;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1485;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [31:0] _RAND_1491;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
  reg [31:0] _RAND_1514;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [31:0] _RAND_1518;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1521;
  reg [31:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1525;
  reg [31:0] _RAND_1526;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [31:0] _RAND_1530;
  reg [31:0] _RAND_1531;
  reg [31:0] _RAND_1532;
  reg [31:0] _RAND_1533;
  reg [31:0] _RAND_1534;
  reg [31:0] _RAND_1535;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1537;
  reg [31:0] _RAND_1538;
  reg [31:0] _RAND_1539;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [31:0] _RAND_1542;
  reg [31:0] _RAND_1543;
`endif // RANDOMIZE_REG_INIT
  wire  adderTreeInst_clock; // @[block_division.scala 223:29]
  wire  adderTreeInst_reset; // @[block_division.scala 223:29]
  wire [5:0] adderTreeInst_io_sign_man_0; // @[block_division.scala 223:29]
  wire [5:0] adderTreeInst_io_sign_man_1; // @[block_division.scala 223:29]
  wire [5:0] adderTreeInst_io_sign_man_2; // @[block_division.scala 223:29]
  wire [5:0] adderTreeInst_io_sign_man_3; // @[block_division.scala 223:29]
  wire [8:0] adderTreeInst_io_exps_0; // @[block_division.scala 223:29]
  wire [8:0] adderTreeInst_io_exps_1; // @[block_division.scala 223:29]
  wire [8:0] adderTreeInst_io_exps_2; // @[block_division.scala 223:29]
  wire [8:0] adderTreeInst_io_exps_3; // @[block_division.scala 223:29]
  wire  adderTreeInst_io_control_signal; // @[block_division.scala 223:29]
  wire  adderTreeInst_io_control_signal2; // @[block_division.scala 223:29]
  wire [13:0] adderTreeInst_io_result_tree; // @[block_division.scala 223:29]
  reg [8:0] exp_output_0; // @[block_division.scala 194:60]
  reg [8:0] exp_output_1; // @[block_division.scala 194:60]
  reg [8:0] exp_output_2; // @[block_division.scala 194:60]
  reg [8:0] exp_output_3; // @[block_division.scala 194:60]
  reg [5:0] acc_0; // @[block_division.scala 195:53]
  reg [5:0] acc_1; // @[block_division.scala 195:53]
  reg [5:0] acc_2; // @[block_division.scala 195:53]
  reg [5:0] acc_3; // @[block_division.scala 195:53]
  wire [8:0] _exp_output_0_T = io_exp_a_0 + io_exp_b_0; // @[block_division.scala 198:34]
  reg [4:0] dotProductRegs__0; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__1; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__2; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__3; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__4; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__5; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__6; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__7; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__8; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__9; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__10; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__11; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__12; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__13; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__14; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__15; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__16; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__17; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__18; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__19; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__20; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__21; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__22; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__23; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__24; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__25; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__26; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__27; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__28; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__29; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__30; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__31; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__32; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__33; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__34; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__35; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__36; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__37; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__38; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__39; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__40; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__41; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__42; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__43; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__44; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__45; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__46; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__47; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__48; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__49; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__50; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__51; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__52; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__53; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__54; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__55; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__56; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__57; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__58; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__59; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__60; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__61; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__62; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs__63; // @[block_division.scala 199:29]
  reg  signs__0; // @[block_division.scala 200:20]
  reg  signs__1; // @[block_division.scala 200:20]
  reg  signs__2; // @[block_division.scala 200:20]
  reg  signs__3; // @[block_division.scala 200:20]
  reg  signs__4; // @[block_division.scala 200:20]
  reg  signs__5; // @[block_division.scala 200:20]
  reg  signs__6; // @[block_division.scala 200:20]
  reg  signs__7; // @[block_division.scala 200:20]
  reg  signs__8; // @[block_division.scala 200:20]
  reg  signs__9; // @[block_division.scala 200:20]
  reg  signs__10; // @[block_division.scala 200:20]
  reg  signs__11; // @[block_division.scala 200:20]
  reg  signs__12; // @[block_division.scala 200:20]
  reg  signs__13; // @[block_division.scala 200:20]
  reg  signs__14; // @[block_division.scala 200:20]
  reg  signs__15; // @[block_division.scala 200:20]
  reg  signs__16; // @[block_division.scala 200:20]
  reg  signs__17; // @[block_division.scala 200:20]
  reg  signs__18; // @[block_division.scala 200:20]
  reg  signs__19; // @[block_division.scala 200:20]
  reg  signs__20; // @[block_division.scala 200:20]
  reg  signs__21; // @[block_division.scala 200:20]
  reg  signs__22; // @[block_division.scala 200:20]
  reg  signs__23; // @[block_division.scala 200:20]
  reg  signs__24; // @[block_division.scala 200:20]
  reg  signs__25; // @[block_division.scala 200:20]
  reg  signs__26; // @[block_division.scala 200:20]
  reg  signs__27; // @[block_division.scala 200:20]
  reg  signs__28; // @[block_division.scala 200:20]
  reg  signs__29; // @[block_division.scala 200:20]
  reg  signs__30; // @[block_division.scala 200:20]
  reg  signs__31; // @[block_division.scala 200:20]
  reg  signs__32; // @[block_division.scala 200:20]
  reg  signs__33; // @[block_division.scala 200:20]
  reg  signs__34; // @[block_division.scala 200:20]
  reg  signs__35; // @[block_division.scala 200:20]
  reg  signs__36; // @[block_division.scala 200:20]
  reg  signs__37; // @[block_division.scala 200:20]
  reg  signs__38; // @[block_division.scala 200:20]
  reg  signs__39; // @[block_division.scala 200:20]
  reg  signs__40; // @[block_division.scala 200:20]
  reg  signs__41; // @[block_division.scala 200:20]
  reg  signs__42; // @[block_division.scala 200:20]
  reg  signs__43; // @[block_division.scala 200:20]
  reg  signs__44; // @[block_division.scala 200:20]
  reg  signs__45; // @[block_division.scala 200:20]
  reg  signs__46; // @[block_division.scala 200:20]
  reg  signs__47; // @[block_division.scala 200:20]
  reg  signs__48; // @[block_division.scala 200:20]
  reg  signs__49; // @[block_division.scala 200:20]
  reg  signs__50; // @[block_division.scala 200:20]
  reg  signs__51; // @[block_division.scala 200:20]
  reg  signs__52; // @[block_division.scala 200:20]
  reg  signs__53; // @[block_division.scala 200:20]
  reg  signs__54; // @[block_division.scala 200:20]
  reg  signs__55; // @[block_division.scala 200:20]
  reg  signs__56; // @[block_division.scala 200:20]
  reg  signs__57; // @[block_division.scala 200:20]
  reg  signs__58; // @[block_division.scala 200:20]
  reg  signs__59; // @[block_division.scala 200:20]
  reg  signs__60; // @[block_division.scala 200:20]
  reg  signs__61; // @[block_division.scala 200:20]
  reg  signs__62; // @[block_division.scala 200:20]
  reg  signs__63; // @[block_division.scala 200:20]
  reg [5:0] two_complement__0; // @[block_division.scala 201:29]
  reg [5:0] two_complement__1; // @[block_division.scala 201:29]
  reg [5:0] two_complement__2; // @[block_division.scala 201:29]
  reg [5:0] two_complement__3; // @[block_division.scala 201:29]
  reg [5:0] two_complement__4; // @[block_division.scala 201:29]
  reg [5:0] two_complement__5; // @[block_division.scala 201:29]
  reg [5:0] two_complement__6; // @[block_division.scala 201:29]
  reg [5:0] two_complement__7; // @[block_division.scala 201:29]
  reg [5:0] two_complement__8; // @[block_division.scala 201:29]
  reg [5:0] two_complement__9; // @[block_division.scala 201:29]
  reg [5:0] two_complement__10; // @[block_division.scala 201:29]
  reg [5:0] two_complement__11; // @[block_division.scala 201:29]
  reg [5:0] two_complement__12; // @[block_division.scala 201:29]
  reg [5:0] two_complement__13; // @[block_division.scala 201:29]
  reg [5:0] two_complement__14; // @[block_division.scala 201:29]
  reg [5:0] two_complement__15; // @[block_division.scala 201:29]
  reg [5:0] two_complement__16; // @[block_division.scala 201:29]
  reg [5:0] two_complement__17; // @[block_division.scala 201:29]
  reg [5:0] two_complement__18; // @[block_division.scala 201:29]
  reg [5:0] two_complement__19; // @[block_division.scala 201:29]
  reg [5:0] two_complement__20; // @[block_division.scala 201:29]
  reg [5:0] two_complement__21; // @[block_division.scala 201:29]
  reg [5:0] two_complement__22; // @[block_division.scala 201:29]
  reg [5:0] two_complement__23; // @[block_division.scala 201:29]
  reg [5:0] two_complement__24; // @[block_division.scala 201:29]
  reg [5:0] two_complement__25; // @[block_division.scala 201:29]
  reg [5:0] two_complement__26; // @[block_division.scala 201:29]
  reg [5:0] two_complement__27; // @[block_division.scala 201:29]
  reg [5:0] two_complement__28; // @[block_division.scala 201:29]
  reg [5:0] two_complement__29; // @[block_division.scala 201:29]
  reg [5:0] two_complement__30; // @[block_division.scala 201:29]
  reg [5:0] two_complement__31; // @[block_division.scala 201:29]
  reg [5:0] two_complement__32; // @[block_division.scala 201:29]
  reg [5:0] two_complement__33; // @[block_division.scala 201:29]
  reg [5:0] two_complement__34; // @[block_division.scala 201:29]
  reg [5:0] two_complement__35; // @[block_division.scala 201:29]
  reg [5:0] two_complement__36; // @[block_division.scala 201:29]
  reg [5:0] two_complement__37; // @[block_division.scala 201:29]
  reg [5:0] two_complement__38; // @[block_division.scala 201:29]
  reg [5:0] two_complement__39; // @[block_division.scala 201:29]
  reg [5:0] two_complement__40; // @[block_division.scala 201:29]
  reg [5:0] two_complement__41; // @[block_division.scala 201:29]
  reg [5:0] two_complement__42; // @[block_division.scala 201:29]
  reg [5:0] two_complement__43; // @[block_division.scala 201:29]
  reg [5:0] two_complement__44; // @[block_division.scala 201:29]
  reg [5:0] two_complement__45; // @[block_division.scala 201:29]
  reg [5:0] two_complement__46; // @[block_division.scala 201:29]
  reg [5:0] two_complement__47; // @[block_division.scala 201:29]
  reg [5:0] two_complement__48; // @[block_division.scala 201:29]
  reg [5:0] two_complement__49; // @[block_division.scala 201:29]
  reg [5:0] two_complement__50; // @[block_division.scala 201:29]
  reg [5:0] two_complement__51; // @[block_division.scala 201:29]
  reg [5:0] two_complement__52; // @[block_division.scala 201:29]
  reg [5:0] two_complement__53; // @[block_division.scala 201:29]
  reg [5:0] two_complement__54; // @[block_division.scala 201:29]
  reg [5:0] two_complement__55; // @[block_division.scala 201:29]
  reg [5:0] two_complement__56; // @[block_division.scala 201:29]
  reg [5:0] two_complement__57; // @[block_division.scala 201:29]
  reg [5:0] two_complement__58; // @[block_division.scala 201:29]
  reg [5:0] two_complement__59; // @[block_division.scala 201:29]
  reg [5:0] two_complement__60; // @[block_division.scala 201:29]
  reg [5:0] two_complement__61; // @[block_division.scala 201:29]
  reg [5:0] two_complement__62; // @[block_division.scala 201:29]
  reg [5:0] two_complement__63; // @[block_division.scala 201:29]
  reg [5:0] two_complement_buffer__0; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__1; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__2; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__3; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__4; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__5; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__6; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__7; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__8; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__9; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__10; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__11; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__12; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__13; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__14; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__15; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__16; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__17; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__18; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__19; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__20; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__21; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__22; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__23; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__24; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__25; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__26; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__27; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__28; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__29; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__30; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__31; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__32; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__33; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__34; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__35; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__36; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__37; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__38; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__39; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__40; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__41; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__42; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__43; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__44; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__45; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__46; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__47; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__48; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__49; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__50; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__51; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__52; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__53; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__54; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__55; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__56; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__57; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__58; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__59; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__60; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__61; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__62; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer__63; // @[block_division.scala 202:36]
  reg [4:0] multiplierReg; // @[block_division.scala 204:34]
  reg  signReg; // @[block_division.scala 205:28]
  wire [9:0] multiplication = multiplierReg * io_man_b_0; // @[block_division.scala 208:42]
  wire [5:0] _dotProductRegs_0_T_1 = 6'h20 - 6'h1; // @[block_division.scala 209:60]
  wire [9:0] _GEN_0 = {{4'd0}, _dotProductRegs_0_T_1}; // @[block_division.scala 209:47]
  wire [9:0] _dotProductRegs_0_T_5 = multiplication > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_0_T_1 = {1'h0,dotProductRegs__0}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_0_T_2 = ~_two_complement_0_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_0_T_4 = _two_complement_0_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_1; // @[block_division.scala 204:34]
  reg  signReg_1; // @[block_division.scala 205:28]
  wire [9:0] multiplication_1 = multiplierReg_1 * io_man_b_1; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_1_T_5 = multiplication_1 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_1; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_1_T_1 = {1'h0,dotProductRegs__1}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_1_T_2 = ~_two_complement_1_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_1_T_4 = _two_complement_1_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_2; // @[block_division.scala 204:34]
  reg  signReg_2; // @[block_division.scala 205:28]
  wire [9:0] multiplication_2 = multiplierReg_2 * io_man_b_2; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_2_T_5 = multiplication_2 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_2; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_2_T_1 = {1'h0,dotProductRegs__2}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_2_T_2 = ~_two_complement_2_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_2_T_4 = _two_complement_2_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_3; // @[block_division.scala 204:34]
  reg  signReg_3; // @[block_division.scala 205:28]
  wire [9:0] multiplication_3 = multiplierReg_3 * io_man_b_3; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_3_T_5 = multiplication_3 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_3; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_3_T_1 = {1'h0,dotProductRegs__3}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_3_T_2 = ~_two_complement_3_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_3_T_4 = _two_complement_3_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_4; // @[block_division.scala 204:34]
  reg  signReg_4; // @[block_division.scala 205:28]
  wire [9:0] multiplication_4 = multiplierReg_4 * io_man_b_4; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_4_T_5 = multiplication_4 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_4; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_4_T_1 = {1'h0,dotProductRegs__4}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_4_T_2 = ~_two_complement_4_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_4_T_4 = _two_complement_4_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_5; // @[block_division.scala 204:34]
  reg  signReg_5; // @[block_division.scala 205:28]
  wire [9:0] multiplication_5 = multiplierReg_5 * io_man_b_5; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_5_T_5 = multiplication_5 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_5; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_5_T_1 = {1'h0,dotProductRegs__5}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_5_T_2 = ~_two_complement_5_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_5_T_4 = _two_complement_5_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_6; // @[block_division.scala 204:34]
  reg  signReg_6; // @[block_division.scala 205:28]
  wire [9:0] multiplication_6 = multiplierReg_6 * io_man_b_6; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_6_T_5 = multiplication_6 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_6; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_6_T_1 = {1'h0,dotProductRegs__6}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_6_T_2 = ~_two_complement_6_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_6_T_4 = _two_complement_6_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_7; // @[block_division.scala 204:34]
  reg  signReg_7; // @[block_division.scala 205:28]
  wire [9:0] multiplication_7 = multiplierReg_7 * io_man_b_7; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_7_T_5 = multiplication_7 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_7; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_7_T_1 = {1'h0,dotProductRegs__7}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_7_T_2 = ~_two_complement_7_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_7_T_4 = _two_complement_7_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_8; // @[block_division.scala 204:34]
  reg  signReg_8; // @[block_division.scala 205:28]
  wire [9:0] multiplication_8 = multiplierReg_8 * io_man_b_8; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_8_T_5 = multiplication_8 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_8; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_8_T_1 = {1'h0,dotProductRegs__8}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_8_T_2 = ~_two_complement_8_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_8_T_4 = _two_complement_8_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_9; // @[block_division.scala 204:34]
  reg  signReg_9; // @[block_division.scala 205:28]
  wire [9:0] multiplication_9 = multiplierReg_9 * io_man_b_9; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_9_T_5 = multiplication_9 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_9; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_9_T_1 = {1'h0,dotProductRegs__9}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_9_T_2 = ~_two_complement_9_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_9_T_4 = _two_complement_9_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_10; // @[block_division.scala 204:34]
  reg  signReg_10; // @[block_division.scala 205:28]
  wire [9:0] multiplication_10 = multiplierReg_10 * io_man_b_10; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_10_T_5 = multiplication_10 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_10; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_10_T_1 = {1'h0,dotProductRegs__10}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_10_T_2 = ~_two_complement_10_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_10_T_4 = _two_complement_10_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_11; // @[block_division.scala 204:34]
  reg  signReg_11; // @[block_division.scala 205:28]
  wire [9:0] multiplication_11 = multiplierReg_11 * io_man_b_11; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_11_T_5 = multiplication_11 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_11; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_11_T_1 = {1'h0,dotProductRegs__11}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_11_T_2 = ~_two_complement_11_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_11_T_4 = _two_complement_11_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_12; // @[block_division.scala 204:34]
  reg  signReg_12; // @[block_division.scala 205:28]
  wire [9:0] multiplication_12 = multiplierReg_12 * io_man_b_12; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_12_T_5 = multiplication_12 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_12; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_12_T_1 = {1'h0,dotProductRegs__12}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_12_T_2 = ~_two_complement_12_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_12_T_4 = _two_complement_12_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_13; // @[block_division.scala 204:34]
  reg  signReg_13; // @[block_division.scala 205:28]
  wire [9:0] multiplication_13 = multiplierReg_13 * io_man_b_13; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_13_T_5 = multiplication_13 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_13; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_13_T_1 = {1'h0,dotProductRegs__13}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_13_T_2 = ~_two_complement_13_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_13_T_4 = _two_complement_13_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_14; // @[block_division.scala 204:34]
  reg  signReg_14; // @[block_division.scala 205:28]
  wire [9:0] multiplication_14 = multiplierReg_14 * io_man_b_14; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_14_T_5 = multiplication_14 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_14; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_14_T_1 = {1'h0,dotProductRegs__14}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_14_T_2 = ~_two_complement_14_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_14_T_4 = _two_complement_14_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_15; // @[block_division.scala 204:34]
  reg  signReg_15; // @[block_division.scala 205:28]
  wire [9:0] multiplication_15 = multiplierReg_15 * io_man_b_15; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_15_T_5 = multiplication_15 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_15; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_15_T_1 = {1'h0,dotProductRegs__15}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_15_T_2 = ~_two_complement_15_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_15_T_4 = _two_complement_15_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_16; // @[block_division.scala 204:34]
  reg  signReg_16; // @[block_division.scala 205:28]
  wire [9:0] multiplication_16 = multiplierReg_16 * io_man_b_16; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_16_T_5 = multiplication_16 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_16; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_16_T_1 = {1'h0,dotProductRegs__16}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_16_T_2 = ~_two_complement_16_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_16_T_4 = _two_complement_16_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_17; // @[block_division.scala 204:34]
  reg  signReg_17; // @[block_division.scala 205:28]
  wire [9:0] multiplication_17 = multiplierReg_17 * io_man_b_17; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_17_T_5 = multiplication_17 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_17; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_17_T_1 = {1'h0,dotProductRegs__17}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_17_T_2 = ~_two_complement_17_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_17_T_4 = _two_complement_17_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_18; // @[block_division.scala 204:34]
  reg  signReg_18; // @[block_division.scala 205:28]
  wire [9:0] multiplication_18 = multiplierReg_18 * io_man_b_18; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_18_T_5 = multiplication_18 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_18; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_18_T_1 = {1'h0,dotProductRegs__18}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_18_T_2 = ~_two_complement_18_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_18_T_4 = _two_complement_18_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_19; // @[block_division.scala 204:34]
  reg  signReg_19; // @[block_division.scala 205:28]
  wire [9:0] multiplication_19 = multiplierReg_19 * io_man_b_19; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_19_T_5 = multiplication_19 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_19; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_19_T_1 = {1'h0,dotProductRegs__19}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_19_T_2 = ~_two_complement_19_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_19_T_4 = _two_complement_19_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_20; // @[block_division.scala 204:34]
  reg  signReg_20; // @[block_division.scala 205:28]
  wire [9:0] multiplication_20 = multiplierReg_20 * io_man_b_20; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_20_T_5 = multiplication_20 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_20; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_20_T_1 = {1'h0,dotProductRegs__20}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_20_T_2 = ~_two_complement_20_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_20_T_4 = _two_complement_20_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_21; // @[block_division.scala 204:34]
  reg  signReg_21; // @[block_division.scala 205:28]
  wire [9:0] multiplication_21 = multiplierReg_21 * io_man_b_21; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_21_T_5 = multiplication_21 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_21; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_21_T_1 = {1'h0,dotProductRegs__21}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_21_T_2 = ~_two_complement_21_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_21_T_4 = _two_complement_21_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_22; // @[block_division.scala 204:34]
  reg  signReg_22; // @[block_division.scala 205:28]
  wire [9:0] multiplication_22 = multiplierReg_22 * io_man_b_22; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_22_T_5 = multiplication_22 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_22; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_22_T_1 = {1'h0,dotProductRegs__22}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_22_T_2 = ~_two_complement_22_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_22_T_4 = _two_complement_22_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_23; // @[block_division.scala 204:34]
  reg  signReg_23; // @[block_division.scala 205:28]
  wire [9:0] multiplication_23 = multiplierReg_23 * io_man_b_23; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_23_T_5 = multiplication_23 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_23; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_23_T_1 = {1'h0,dotProductRegs__23}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_23_T_2 = ~_two_complement_23_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_23_T_4 = _two_complement_23_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_24; // @[block_division.scala 204:34]
  reg  signReg_24; // @[block_division.scala 205:28]
  wire [9:0] multiplication_24 = multiplierReg_24 * io_man_b_24; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_24_T_5 = multiplication_24 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_24; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_24_T_1 = {1'h0,dotProductRegs__24}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_24_T_2 = ~_two_complement_24_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_24_T_4 = _two_complement_24_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_25; // @[block_division.scala 204:34]
  reg  signReg_25; // @[block_division.scala 205:28]
  wire [9:0] multiplication_25 = multiplierReg_25 * io_man_b_25; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_25_T_5 = multiplication_25 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_25; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_25_T_1 = {1'h0,dotProductRegs__25}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_25_T_2 = ~_two_complement_25_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_25_T_4 = _two_complement_25_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_26; // @[block_division.scala 204:34]
  reg  signReg_26; // @[block_division.scala 205:28]
  wire [9:0] multiplication_26 = multiplierReg_26 * io_man_b_26; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_26_T_5 = multiplication_26 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_26; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_26_T_1 = {1'h0,dotProductRegs__26}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_26_T_2 = ~_two_complement_26_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_26_T_4 = _two_complement_26_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_27; // @[block_division.scala 204:34]
  reg  signReg_27; // @[block_division.scala 205:28]
  wire [9:0] multiplication_27 = multiplierReg_27 * io_man_b_27; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_27_T_5 = multiplication_27 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_27; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_27_T_1 = {1'h0,dotProductRegs__27}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_27_T_2 = ~_two_complement_27_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_27_T_4 = _two_complement_27_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_28; // @[block_division.scala 204:34]
  reg  signReg_28; // @[block_division.scala 205:28]
  wire [9:0] multiplication_28 = multiplierReg_28 * io_man_b_28; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_28_T_5 = multiplication_28 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_28; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_28_T_1 = {1'h0,dotProductRegs__28}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_28_T_2 = ~_two_complement_28_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_28_T_4 = _two_complement_28_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_29; // @[block_division.scala 204:34]
  reg  signReg_29; // @[block_division.scala 205:28]
  wire [9:0] multiplication_29 = multiplierReg_29 * io_man_b_29; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_29_T_5 = multiplication_29 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_29; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_29_T_1 = {1'h0,dotProductRegs__29}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_29_T_2 = ~_two_complement_29_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_29_T_4 = _two_complement_29_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_30; // @[block_division.scala 204:34]
  reg  signReg_30; // @[block_division.scala 205:28]
  wire [9:0] multiplication_30 = multiplierReg_30 * io_man_b_30; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_30_T_5 = multiplication_30 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_30; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_30_T_1 = {1'h0,dotProductRegs__30}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_30_T_2 = ~_two_complement_30_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_30_T_4 = _two_complement_30_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_31; // @[block_division.scala 204:34]
  reg  signReg_31; // @[block_division.scala 205:28]
  wire [9:0] multiplication_31 = multiplierReg_31 * io_man_b_31; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_31_T_5 = multiplication_31 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_31; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_31_T_1 = {1'h0,dotProductRegs__31}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_31_T_2 = ~_two_complement_31_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_31_T_4 = _two_complement_31_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_32; // @[block_division.scala 204:34]
  reg  signReg_32; // @[block_division.scala 205:28]
  wire [9:0] multiplication_32 = multiplierReg_32 * io_man_b_32; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_32_T_5 = multiplication_32 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_32; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_32_T_1 = {1'h0,dotProductRegs__32}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_32_T_2 = ~_two_complement_32_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_32_T_4 = _two_complement_32_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_33; // @[block_division.scala 204:34]
  reg  signReg_33; // @[block_division.scala 205:28]
  wire [9:0] multiplication_33 = multiplierReg_33 * io_man_b_33; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_33_T_5 = multiplication_33 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_33; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_33_T_1 = {1'h0,dotProductRegs__33}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_33_T_2 = ~_two_complement_33_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_33_T_4 = _two_complement_33_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_34; // @[block_division.scala 204:34]
  reg  signReg_34; // @[block_division.scala 205:28]
  wire [9:0] multiplication_34 = multiplierReg_34 * io_man_b_34; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_34_T_5 = multiplication_34 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_34; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_34_T_1 = {1'h0,dotProductRegs__34}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_34_T_2 = ~_two_complement_34_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_34_T_4 = _two_complement_34_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_35; // @[block_division.scala 204:34]
  reg  signReg_35; // @[block_division.scala 205:28]
  wire [9:0] multiplication_35 = multiplierReg_35 * io_man_b_35; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_35_T_5 = multiplication_35 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_35; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_35_T_1 = {1'h0,dotProductRegs__35}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_35_T_2 = ~_two_complement_35_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_35_T_4 = _two_complement_35_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_36; // @[block_division.scala 204:34]
  reg  signReg_36; // @[block_division.scala 205:28]
  wire [9:0] multiplication_36 = multiplierReg_36 * io_man_b_36; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_36_T_5 = multiplication_36 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_36; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_36_T_1 = {1'h0,dotProductRegs__36}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_36_T_2 = ~_two_complement_36_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_36_T_4 = _two_complement_36_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_37; // @[block_division.scala 204:34]
  reg  signReg_37; // @[block_division.scala 205:28]
  wire [9:0] multiplication_37 = multiplierReg_37 * io_man_b_37; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_37_T_5 = multiplication_37 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_37; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_37_T_1 = {1'h0,dotProductRegs__37}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_37_T_2 = ~_two_complement_37_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_37_T_4 = _two_complement_37_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_38; // @[block_division.scala 204:34]
  reg  signReg_38; // @[block_division.scala 205:28]
  wire [9:0] multiplication_38 = multiplierReg_38 * io_man_b_38; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_38_T_5 = multiplication_38 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_38; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_38_T_1 = {1'h0,dotProductRegs__38}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_38_T_2 = ~_two_complement_38_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_38_T_4 = _two_complement_38_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_39; // @[block_division.scala 204:34]
  reg  signReg_39; // @[block_division.scala 205:28]
  wire [9:0] multiplication_39 = multiplierReg_39 * io_man_b_39; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_39_T_5 = multiplication_39 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_39; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_39_T_1 = {1'h0,dotProductRegs__39}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_39_T_2 = ~_two_complement_39_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_39_T_4 = _two_complement_39_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_40; // @[block_division.scala 204:34]
  reg  signReg_40; // @[block_division.scala 205:28]
  wire [9:0] multiplication_40 = multiplierReg_40 * io_man_b_40; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_40_T_5 = multiplication_40 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_40; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_40_T_1 = {1'h0,dotProductRegs__40}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_40_T_2 = ~_two_complement_40_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_40_T_4 = _two_complement_40_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_41; // @[block_division.scala 204:34]
  reg  signReg_41; // @[block_division.scala 205:28]
  wire [9:0] multiplication_41 = multiplierReg_41 * io_man_b_41; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_41_T_5 = multiplication_41 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_41; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_41_T_1 = {1'h0,dotProductRegs__41}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_41_T_2 = ~_two_complement_41_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_41_T_4 = _two_complement_41_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_42; // @[block_division.scala 204:34]
  reg  signReg_42; // @[block_division.scala 205:28]
  wire [9:0] multiplication_42 = multiplierReg_42 * io_man_b_42; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_42_T_5 = multiplication_42 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_42; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_42_T_1 = {1'h0,dotProductRegs__42}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_42_T_2 = ~_two_complement_42_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_42_T_4 = _two_complement_42_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_43; // @[block_division.scala 204:34]
  reg  signReg_43; // @[block_division.scala 205:28]
  wire [9:0] multiplication_43 = multiplierReg_43 * io_man_b_43; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_43_T_5 = multiplication_43 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_43; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_43_T_1 = {1'h0,dotProductRegs__43}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_43_T_2 = ~_two_complement_43_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_43_T_4 = _two_complement_43_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_44; // @[block_division.scala 204:34]
  reg  signReg_44; // @[block_division.scala 205:28]
  wire [9:0] multiplication_44 = multiplierReg_44 * io_man_b_44; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_44_T_5 = multiplication_44 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_44; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_44_T_1 = {1'h0,dotProductRegs__44}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_44_T_2 = ~_two_complement_44_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_44_T_4 = _two_complement_44_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_45; // @[block_division.scala 204:34]
  reg  signReg_45; // @[block_division.scala 205:28]
  wire [9:0] multiplication_45 = multiplierReg_45 * io_man_b_45; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_45_T_5 = multiplication_45 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_45; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_45_T_1 = {1'h0,dotProductRegs__45}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_45_T_2 = ~_two_complement_45_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_45_T_4 = _two_complement_45_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_46; // @[block_division.scala 204:34]
  reg  signReg_46; // @[block_division.scala 205:28]
  wire [9:0] multiplication_46 = multiplierReg_46 * io_man_b_46; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_46_T_5 = multiplication_46 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_46; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_46_T_1 = {1'h0,dotProductRegs__46}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_46_T_2 = ~_two_complement_46_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_46_T_4 = _two_complement_46_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_47; // @[block_division.scala 204:34]
  reg  signReg_47; // @[block_division.scala 205:28]
  wire [9:0] multiplication_47 = multiplierReg_47 * io_man_b_47; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_47_T_5 = multiplication_47 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_47; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_47_T_1 = {1'h0,dotProductRegs__47}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_47_T_2 = ~_two_complement_47_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_47_T_4 = _two_complement_47_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_48; // @[block_division.scala 204:34]
  reg  signReg_48; // @[block_division.scala 205:28]
  wire [9:0] multiplication_48 = multiplierReg_48 * io_man_b_48; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_48_T_5 = multiplication_48 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_48; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_48_T_1 = {1'h0,dotProductRegs__48}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_48_T_2 = ~_two_complement_48_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_48_T_4 = _two_complement_48_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_49; // @[block_division.scala 204:34]
  reg  signReg_49; // @[block_division.scala 205:28]
  wire [9:0] multiplication_49 = multiplierReg_49 * io_man_b_49; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_49_T_5 = multiplication_49 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_49; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_49_T_1 = {1'h0,dotProductRegs__49}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_49_T_2 = ~_two_complement_49_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_49_T_4 = _two_complement_49_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_50; // @[block_division.scala 204:34]
  reg  signReg_50; // @[block_division.scala 205:28]
  wire [9:0] multiplication_50 = multiplierReg_50 * io_man_b_50; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_50_T_5 = multiplication_50 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_50; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_50_T_1 = {1'h0,dotProductRegs__50}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_50_T_2 = ~_two_complement_50_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_50_T_4 = _two_complement_50_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_51; // @[block_division.scala 204:34]
  reg  signReg_51; // @[block_division.scala 205:28]
  wire [9:0] multiplication_51 = multiplierReg_51 * io_man_b_51; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_51_T_5 = multiplication_51 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_51; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_51_T_1 = {1'h0,dotProductRegs__51}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_51_T_2 = ~_two_complement_51_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_51_T_4 = _two_complement_51_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_52; // @[block_division.scala 204:34]
  reg  signReg_52; // @[block_division.scala 205:28]
  wire [9:0] multiplication_52 = multiplierReg_52 * io_man_b_52; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_52_T_5 = multiplication_52 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_52; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_52_T_1 = {1'h0,dotProductRegs__52}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_52_T_2 = ~_two_complement_52_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_52_T_4 = _two_complement_52_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_53; // @[block_division.scala 204:34]
  reg  signReg_53; // @[block_division.scala 205:28]
  wire [9:0] multiplication_53 = multiplierReg_53 * io_man_b_53; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_53_T_5 = multiplication_53 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_53; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_53_T_1 = {1'h0,dotProductRegs__53}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_53_T_2 = ~_two_complement_53_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_53_T_4 = _two_complement_53_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_54; // @[block_division.scala 204:34]
  reg  signReg_54; // @[block_division.scala 205:28]
  wire [9:0] multiplication_54 = multiplierReg_54 * io_man_b_54; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_54_T_5 = multiplication_54 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_54; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_54_T_1 = {1'h0,dotProductRegs__54}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_54_T_2 = ~_two_complement_54_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_54_T_4 = _two_complement_54_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_55; // @[block_division.scala 204:34]
  reg  signReg_55; // @[block_division.scala 205:28]
  wire [9:0] multiplication_55 = multiplierReg_55 * io_man_b_55; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_55_T_5 = multiplication_55 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_55; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_55_T_1 = {1'h0,dotProductRegs__55}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_55_T_2 = ~_two_complement_55_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_55_T_4 = _two_complement_55_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_56; // @[block_division.scala 204:34]
  reg  signReg_56; // @[block_division.scala 205:28]
  wire [9:0] multiplication_56 = multiplierReg_56 * io_man_b_56; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_56_T_5 = multiplication_56 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_56; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_56_T_1 = {1'h0,dotProductRegs__56}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_56_T_2 = ~_two_complement_56_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_56_T_4 = _two_complement_56_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_57; // @[block_division.scala 204:34]
  reg  signReg_57; // @[block_division.scala 205:28]
  wire [9:0] multiplication_57 = multiplierReg_57 * io_man_b_57; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_57_T_5 = multiplication_57 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_57; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_57_T_1 = {1'h0,dotProductRegs__57}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_57_T_2 = ~_two_complement_57_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_57_T_4 = _two_complement_57_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_58; // @[block_division.scala 204:34]
  reg  signReg_58; // @[block_division.scala 205:28]
  wire [9:0] multiplication_58 = multiplierReg_58 * io_man_b_58; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_58_T_5 = multiplication_58 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_58; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_58_T_1 = {1'h0,dotProductRegs__58}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_58_T_2 = ~_two_complement_58_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_58_T_4 = _two_complement_58_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_59; // @[block_division.scala 204:34]
  reg  signReg_59; // @[block_division.scala 205:28]
  wire [9:0] multiplication_59 = multiplierReg_59 * io_man_b_59; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_59_T_5 = multiplication_59 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_59; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_59_T_1 = {1'h0,dotProductRegs__59}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_59_T_2 = ~_two_complement_59_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_59_T_4 = _two_complement_59_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_60; // @[block_division.scala 204:34]
  reg  signReg_60; // @[block_division.scala 205:28]
  wire [9:0] multiplication_60 = multiplierReg_60 * io_man_b_60; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_60_T_5 = multiplication_60 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_60; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_60_T_1 = {1'h0,dotProductRegs__60}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_60_T_2 = ~_two_complement_60_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_60_T_4 = _two_complement_60_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_61; // @[block_division.scala 204:34]
  reg  signReg_61; // @[block_division.scala 205:28]
  wire [9:0] multiplication_61 = multiplierReg_61 * io_man_b_61; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_61_T_5 = multiplication_61 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_61; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_61_T_1 = {1'h0,dotProductRegs__61}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_61_T_2 = ~_two_complement_61_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_61_T_4 = _two_complement_61_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_62; // @[block_division.scala 204:34]
  reg  signReg_62; // @[block_division.scala 205:28]
  wire [9:0] multiplication_62 = multiplierReg_62 * io_man_b_62; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_62_T_5 = multiplication_62 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_62; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_62_T_1 = {1'h0,dotProductRegs__62}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_62_T_2 = ~_two_complement_62_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_62_T_4 = _two_complement_62_T_2 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_63; // @[block_division.scala 204:34]
  reg  signReg_63; // @[block_division.scala 205:28]
  wire [9:0] multiplication_63 = multiplierReg_63 * io_man_b_63; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_63_T_5 = multiplication_63 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_63; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_63_T_1 = {1'h0,dotProductRegs__63}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_63_T_2 = ~_two_complement_63_T_1; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_63_T_4 = _two_complement_63_T_2 + 6'h1; // @[block_division.scala 213:38]
  wire [6:0] _sum_T = $signed(two_complement_buffer__0) + $signed(two_complement_buffer__1); // @[block_division.scala 218:46]
  wire [6:0] _GEN_64 = {{1{two_complement_buffer__2[5]}},two_complement_buffer__2}; // @[block_division.scala 218:46]
  wire [7:0] _sum_T_1 = $signed(_sum_T) + $signed(_GEN_64); // @[block_division.scala 218:46]
  wire [7:0] _GEN_65 = {{2{two_complement_buffer__3[5]}},two_complement_buffer__3}; // @[block_division.scala 218:46]
  wire [8:0] _sum_T_2 = $signed(_sum_T_1) + $signed(_GEN_65); // @[block_division.scala 218:46]
  wire [8:0] _GEN_66 = {{3{two_complement_buffer__4[5]}},two_complement_buffer__4}; // @[block_division.scala 218:46]
  wire [9:0] _sum_T_3 = $signed(_sum_T_2) + $signed(_GEN_66); // @[block_division.scala 218:46]
  wire [9:0] _GEN_67 = {{4{two_complement_buffer__5[5]}},two_complement_buffer__5}; // @[block_division.scala 218:46]
  wire [10:0] _sum_T_4 = $signed(_sum_T_3) + $signed(_GEN_67); // @[block_division.scala 218:46]
  wire [10:0] _GEN_68 = {{5{two_complement_buffer__6[5]}},two_complement_buffer__6}; // @[block_division.scala 218:46]
  wire [11:0] _sum_T_5 = $signed(_sum_T_4) + $signed(_GEN_68); // @[block_division.scala 218:46]
  wire [11:0] _GEN_69 = {{6{two_complement_buffer__7[5]}},two_complement_buffer__7}; // @[block_division.scala 218:46]
  wire [12:0] _sum_T_6 = $signed(_sum_T_5) + $signed(_GEN_69); // @[block_division.scala 218:46]
  wire [12:0] _GEN_70 = {{7{two_complement_buffer__8[5]}},two_complement_buffer__8}; // @[block_division.scala 218:46]
  wire [13:0] _sum_T_7 = $signed(_sum_T_6) + $signed(_GEN_70); // @[block_division.scala 218:46]
  wire [13:0] _GEN_71 = {{8{two_complement_buffer__9[5]}},two_complement_buffer__9}; // @[block_division.scala 218:46]
  wire [14:0] _sum_T_8 = $signed(_sum_T_7) + $signed(_GEN_71); // @[block_division.scala 218:46]
  wire [14:0] _GEN_72 = {{9{two_complement_buffer__10[5]}},two_complement_buffer__10}; // @[block_division.scala 218:46]
  wire [15:0] _sum_T_9 = $signed(_sum_T_8) + $signed(_GEN_72); // @[block_division.scala 218:46]
  wire [15:0] _GEN_73 = {{10{two_complement_buffer__11[5]}},two_complement_buffer__11}; // @[block_division.scala 218:46]
  wire [16:0] _sum_T_10 = $signed(_sum_T_9) + $signed(_GEN_73); // @[block_division.scala 218:46]
  wire [16:0] _GEN_74 = {{11{two_complement_buffer__12[5]}},two_complement_buffer__12}; // @[block_division.scala 218:46]
  wire [17:0] _sum_T_11 = $signed(_sum_T_10) + $signed(_GEN_74); // @[block_division.scala 218:46]
  wire [17:0] _GEN_75 = {{12{two_complement_buffer__13[5]}},two_complement_buffer__13}; // @[block_division.scala 218:46]
  wire [18:0] _sum_T_12 = $signed(_sum_T_11) + $signed(_GEN_75); // @[block_division.scala 218:46]
  wire [18:0] _GEN_76 = {{13{two_complement_buffer__14[5]}},two_complement_buffer__14}; // @[block_division.scala 218:46]
  wire [19:0] _sum_T_13 = $signed(_sum_T_12) + $signed(_GEN_76); // @[block_division.scala 218:46]
  wire [19:0] _GEN_77 = {{14{two_complement_buffer__15[5]}},two_complement_buffer__15}; // @[block_division.scala 218:46]
  wire [20:0] _sum_T_14 = $signed(_sum_T_13) + $signed(_GEN_77); // @[block_division.scala 218:46]
  wire [20:0] _GEN_78 = {{15{two_complement_buffer__16[5]}},two_complement_buffer__16}; // @[block_division.scala 218:46]
  wire [21:0] _sum_T_15 = $signed(_sum_T_14) + $signed(_GEN_78); // @[block_division.scala 218:46]
  wire [21:0] _GEN_79 = {{16{two_complement_buffer__17[5]}},two_complement_buffer__17}; // @[block_division.scala 218:46]
  wire [22:0] _sum_T_16 = $signed(_sum_T_15) + $signed(_GEN_79); // @[block_division.scala 218:46]
  wire [22:0] _GEN_80 = {{17{two_complement_buffer__18[5]}},two_complement_buffer__18}; // @[block_division.scala 218:46]
  wire [23:0] _sum_T_17 = $signed(_sum_T_16) + $signed(_GEN_80); // @[block_division.scala 218:46]
  wire [23:0] _GEN_81 = {{18{two_complement_buffer__19[5]}},two_complement_buffer__19}; // @[block_division.scala 218:46]
  wire [24:0] _sum_T_18 = $signed(_sum_T_17) + $signed(_GEN_81); // @[block_division.scala 218:46]
  wire [24:0] _GEN_82 = {{19{two_complement_buffer__20[5]}},two_complement_buffer__20}; // @[block_division.scala 218:46]
  wire [25:0] _sum_T_19 = $signed(_sum_T_18) + $signed(_GEN_82); // @[block_division.scala 218:46]
  wire [25:0] _GEN_83 = {{20{two_complement_buffer__21[5]}},two_complement_buffer__21}; // @[block_division.scala 218:46]
  wire [26:0] _sum_T_20 = $signed(_sum_T_19) + $signed(_GEN_83); // @[block_division.scala 218:46]
  wire [26:0] _GEN_84 = {{21{two_complement_buffer__22[5]}},two_complement_buffer__22}; // @[block_division.scala 218:46]
  wire [27:0] _sum_T_21 = $signed(_sum_T_20) + $signed(_GEN_84); // @[block_division.scala 218:46]
  wire [27:0] _GEN_85 = {{22{two_complement_buffer__23[5]}},two_complement_buffer__23}; // @[block_division.scala 218:46]
  wire [28:0] _sum_T_22 = $signed(_sum_T_21) + $signed(_GEN_85); // @[block_division.scala 218:46]
  wire [28:0] _GEN_86 = {{23{two_complement_buffer__24[5]}},two_complement_buffer__24}; // @[block_division.scala 218:46]
  wire [29:0] _sum_T_23 = $signed(_sum_T_22) + $signed(_GEN_86); // @[block_division.scala 218:46]
  wire [29:0] _GEN_87 = {{24{two_complement_buffer__25[5]}},two_complement_buffer__25}; // @[block_division.scala 218:46]
  wire [30:0] _sum_T_24 = $signed(_sum_T_23) + $signed(_GEN_87); // @[block_division.scala 218:46]
  wire [30:0] _GEN_88 = {{25{two_complement_buffer__26[5]}},two_complement_buffer__26}; // @[block_division.scala 218:46]
  wire [31:0] _sum_T_25 = $signed(_sum_T_24) + $signed(_GEN_88); // @[block_division.scala 218:46]
  wire [31:0] _GEN_89 = {{26{two_complement_buffer__27[5]}},two_complement_buffer__27}; // @[block_division.scala 218:46]
  wire [32:0] _sum_T_26 = $signed(_sum_T_25) + $signed(_GEN_89); // @[block_division.scala 218:46]
  wire [32:0] _GEN_90 = {{27{two_complement_buffer__28[5]}},two_complement_buffer__28}; // @[block_division.scala 218:46]
  wire [33:0] _sum_T_27 = $signed(_sum_T_26) + $signed(_GEN_90); // @[block_division.scala 218:46]
  wire [33:0] _GEN_91 = {{28{two_complement_buffer__29[5]}},two_complement_buffer__29}; // @[block_division.scala 218:46]
  wire [34:0] _sum_T_28 = $signed(_sum_T_27) + $signed(_GEN_91); // @[block_division.scala 218:46]
  wire [34:0] _GEN_92 = {{29{two_complement_buffer__30[5]}},two_complement_buffer__30}; // @[block_division.scala 218:46]
  wire [35:0] _sum_T_29 = $signed(_sum_T_28) + $signed(_GEN_92); // @[block_division.scala 218:46]
  wire [35:0] _GEN_93 = {{30{two_complement_buffer__31[5]}},two_complement_buffer__31}; // @[block_division.scala 218:46]
  wire [36:0] _sum_T_30 = $signed(_sum_T_29) + $signed(_GEN_93); // @[block_division.scala 218:46]
  wire [36:0] _GEN_94 = {{31{two_complement_buffer__32[5]}},two_complement_buffer__32}; // @[block_division.scala 218:46]
  wire [37:0] _sum_T_31 = $signed(_sum_T_30) + $signed(_GEN_94); // @[block_division.scala 218:46]
  wire [37:0] _GEN_95 = {{32{two_complement_buffer__33[5]}},two_complement_buffer__33}; // @[block_division.scala 218:46]
  wire [38:0] _sum_T_32 = $signed(_sum_T_31) + $signed(_GEN_95); // @[block_division.scala 218:46]
  wire [38:0] _GEN_96 = {{33{two_complement_buffer__34[5]}},two_complement_buffer__34}; // @[block_division.scala 218:46]
  wire [39:0] _sum_T_33 = $signed(_sum_T_32) + $signed(_GEN_96); // @[block_division.scala 218:46]
  wire [39:0] _GEN_97 = {{34{two_complement_buffer__35[5]}},two_complement_buffer__35}; // @[block_division.scala 218:46]
  wire [40:0] _sum_T_34 = $signed(_sum_T_33) + $signed(_GEN_97); // @[block_division.scala 218:46]
  wire [40:0] _GEN_98 = {{35{two_complement_buffer__36[5]}},two_complement_buffer__36}; // @[block_division.scala 218:46]
  wire [41:0] _sum_T_35 = $signed(_sum_T_34) + $signed(_GEN_98); // @[block_division.scala 218:46]
  wire [41:0] _GEN_99 = {{36{two_complement_buffer__37[5]}},two_complement_buffer__37}; // @[block_division.scala 218:46]
  wire [42:0] _sum_T_36 = $signed(_sum_T_35) + $signed(_GEN_99); // @[block_division.scala 218:46]
  wire [42:0] _GEN_100 = {{37{two_complement_buffer__38[5]}},two_complement_buffer__38}; // @[block_division.scala 218:46]
  wire [43:0] _sum_T_37 = $signed(_sum_T_36) + $signed(_GEN_100); // @[block_division.scala 218:46]
  wire [43:0] _GEN_101 = {{38{two_complement_buffer__39[5]}},two_complement_buffer__39}; // @[block_division.scala 218:46]
  wire [44:0] _sum_T_38 = $signed(_sum_T_37) + $signed(_GEN_101); // @[block_division.scala 218:46]
  wire [44:0] _GEN_102 = {{39{two_complement_buffer__40[5]}},two_complement_buffer__40}; // @[block_division.scala 218:46]
  wire [45:0] _sum_T_39 = $signed(_sum_T_38) + $signed(_GEN_102); // @[block_division.scala 218:46]
  wire [45:0] _GEN_103 = {{40{two_complement_buffer__41[5]}},two_complement_buffer__41}; // @[block_division.scala 218:46]
  wire [46:0] _sum_T_40 = $signed(_sum_T_39) + $signed(_GEN_103); // @[block_division.scala 218:46]
  wire [46:0] _GEN_104 = {{41{two_complement_buffer__42[5]}},two_complement_buffer__42}; // @[block_division.scala 218:46]
  wire [47:0] _sum_T_41 = $signed(_sum_T_40) + $signed(_GEN_104); // @[block_division.scala 218:46]
  wire [47:0] _GEN_105 = {{42{two_complement_buffer__43[5]}},two_complement_buffer__43}; // @[block_division.scala 218:46]
  wire [48:0] _sum_T_42 = $signed(_sum_T_41) + $signed(_GEN_105); // @[block_division.scala 218:46]
  wire [48:0] _GEN_106 = {{43{two_complement_buffer__44[5]}},two_complement_buffer__44}; // @[block_division.scala 218:46]
  wire [49:0] _sum_T_43 = $signed(_sum_T_42) + $signed(_GEN_106); // @[block_division.scala 218:46]
  wire [49:0] _GEN_107 = {{44{two_complement_buffer__45[5]}},two_complement_buffer__45}; // @[block_division.scala 218:46]
  wire [50:0] _sum_T_44 = $signed(_sum_T_43) + $signed(_GEN_107); // @[block_division.scala 218:46]
  wire [50:0] _GEN_108 = {{45{two_complement_buffer__46[5]}},two_complement_buffer__46}; // @[block_division.scala 218:46]
  wire [51:0] _sum_T_45 = $signed(_sum_T_44) + $signed(_GEN_108); // @[block_division.scala 218:46]
  wire [51:0] _GEN_109 = {{46{two_complement_buffer__47[5]}},two_complement_buffer__47}; // @[block_division.scala 218:46]
  wire [52:0] _sum_T_46 = $signed(_sum_T_45) + $signed(_GEN_109); // @[block_division.scala 218:46]
  wire [52:0] _GEN_110 = {{47{two_complement_buffer__48[5]}},two_complement_buffer__48}; // @[block_division.scala 218:46]
  wire [53:0] _sum_T_47 = $signed(_sum_T_46) + $signed(_GEN_110); // @[block_division.scala 218:46]
  wire [53:0] _GEN_111 = {{48{two_complement_buffer__49[5]}},two_complement_buffer__49}; // @[block_division.scala 218:46]
  wire [54:0] _sum_T_48 = $signed(_sum_T_47) + $signed(_GEN_111); // @[block_division.scala 218:46]
  wire [54:0] _GEN_112 = {{49{two_complement_buffer__50[5]}},two_complement_buffer__50}; // @[block_division.scala 218:46]
  wire [55:0] _sum_T_49 = $signed(_sum_T_48) + $signed(_GEN_112); // @[block_division.scala 218:46]
  wire [55:0] _GEN_113 = {{50{two_complement_buffer__51[5]}},two_complement_buffer__51}; // @[block_division.scala 218:46]
  wire [56:0] _sum_T_50 = $signed(_sum_T_49) + $signed(_GEN_113); // @[block_division.scala 218:46]
  wire [56:0] _GEN_114 = {{51{two_complement_buffer__52[5]}},two_complement_buffer__52}; // @[block_division.scala 218:46]
  wire [57:0] _sum_T_51 = $signed(_sum_T_50) + $signed(_GEN_114); // @[block_division.scala 218:46]
  wire [57:0] _GEN_115 = {{52{two_complement_buffer__53[5]}},two_complement_buffer__53}; // @[block_division.scala 218:46]
  wire [58:0] _sum_T_52 = $signed(_sum_T_51) + $signed(_GEN_115); // @[block_division.scala 218:46]
  wire [58:0] _GEN_116 = {{53{two_complement_buffer__54[5]}},two_complement_buffer__54}; // @[block_division.scala 218:46]
  wire [59:0] _sum_T_53 = $signed(_sum_T_52) + $signed(_GEN_116); // @[block_division.scala 218:46]
  wire [59:0] _GEN_117 = {{54{two_complement_buffer__55[5]}},two_complement_buffer__55}; // @[block_division.scala 218:46]
  wire [60:0] _sum_T_54 = $signed(_sum_T_53) + $signed(_GEN_117); // @[block_division.scala 218:46]
  wire [60:0] _GEN_118 = {{55{two_complement_buffer__56[5]}},two_complement_buffer__56}; // @[block_division.scala 218:46]
  wire [61:0] _sum_T_55 = $signed(_sum_T_54) + $signed(_GEN_118); // @[block_division.scala 218:46]
  wire [61:0] _GEN_119 = {{56{two_complement_buffer__57[5]}},two_complement_buffer__57}; // @[block_division.scala 218:46]
  wire [62:0] _sum_T_56 = $signed(_sum_T_55) + $signed(_GEN_119); // @[block_division.scala 218:46]
  wire [62:0] _GEN_120 = {{57{two_complement_buffer__58[5]}},two_complement_buffer__58}; // @[block_division.scala 218:46]
  wire [63:0] _sum_T_57 = $signed(_sum_T_56) + $signed(_GEN_120); // @[block_division.scala 218:46]
  wire [63:0] _GEN_121 = {{58{two_complement_buffer__59[5]}},two_complement_buffer__59}; // @[block_division.scala 218:46]
  wire [64:0] _sum_T_58 = $signed(_sum_T_57) + $signed(_GEN_121); // @[block_division.scala 218:46]
  wire [64:0] _GEN_122 = {{59{two_complement_buffer__60[5]}},two_complement_buffer__60}; // @[block_division.scala 218:46]
  wire [65:0] _sum_T_59 = $signed(_sum_T_58) + $signed(_GEN_122); // @[block_division.scala 218:46]
  wire [65:0] _GEN_123 = {{60{two_complement_buffer__61[5]}},two_complement_buffer__61}; // @[block_division.scala 218:46]
  wire [66:0] _sum_T_60 = $signed(_sum_T_59) + $signed(_GEN_123); // @[block_division.scala 218:46]
  wire [66:0] _GEN_124 = {{61{two_complement_buffer__62[5]}},two_complement_buffer__62}; // @[block_division.scala 218:46]
  wire [67:0] _sum_T_61 = $signed(_sum_T_60) + $signed(_GEN_124); // @[block_division.scala 218:46]
  wire [67:0] _GEN_125 = {{62{two_complement_buffer__63[5]}},two_complement_buffer__63}; // @[block_division.scala 218:46]
  wire [68:0] sum = $signed(_sum_T_61) + $signed(_GEN_125); // @[block_division.scala 218:46]
  wire [67:0] _acc_0_T_3 = ~sum[67:0]; // @[block_division.scala 219:57]
  wire [67:0] _acc_0_T_5 = _acc_0_T_3 + 68'h1; // @[block_division.scala 219:86]
  wire [67:0] _GEN_126 = {{62'd0}, _dotProductRegs_0_T_1}; // @[block_division.scala 219:93]
  wire [5:0] _acc_0_T_11 = ~_dotProductRegs_0_T_1; // @[block_division.scala 219:114]
  wire [5:0] _acc_0_T_13 = _acc_0_T_11 + 6'h1; // @[block_division.scala 219:135]
  wire [68:0] _acc_0_T_14 = $signed(_sum_T_61) + $signed(_GEN_125); // @[block_division.scala 219:145]
  wire [68:0] _acc_0_T_15 = _acc_0_T_5 > _GEN_126 ? {{63'd0}, _acc_0_T_13} : _acc_0_T_14; // @[block_division.scala 219:55]
  wire [68:0] _acc_0_T_23 = sum[67:0] > _GEN_126 ? {{63'd0}, _dotProductRegs_0_T_1} : _acc_0_T_14; // @[block_division.scala 220:6]
  wire [68:0] _acc_0_T_24 = sum[68] ? _acc_0_T_15 : _acc_0_T_23; // @[block_division.scala 219:18]
  wire [8:0] _exp_output_1_T = io_exp_a_1 + io_exp_b_1; // @[block_division.scala 198:34]
  reg [4:0] dotProductRegs_1_0; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_1; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_2; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_3; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_4; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_5; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_6; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_7; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_8; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_9; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_10; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_11; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_12; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_13; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_14; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_15; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_16; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_17; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_18; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_19; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_20; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_21; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_22; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_23; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_24; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_25; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_26; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_27; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_28; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_29; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_30; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_31; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_32; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_33; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_34; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_35; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_36; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_37; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_38; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_39; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_40; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_41; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_42; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_43; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_44; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_45; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_46; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_47; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_48; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_49; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_50; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_51; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_52; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_53; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_54; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_55; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_56; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_57; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_58; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_59; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_60; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_61; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_62; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_1_63; // @[block_division.scala 199:29]
  reg  signs_1_0; // @[block_division.scala 200:20]
  reg  signs_1_1; // @[block_division.scala 200:20]
  reg  signs_1_2; // @[block_division.scala 200:20]
  reg  signs_1_3; // @[block_division.scala 200:20]
  reg  signs_1_4; // @[block_division.scala 200:20]
  reg  signs_1_5; // @[block_division.scala 200:20]
  reg  signs_1_6; // @[block_division.scala 200:20]
  reg  signs_1_7; // @[block_division.scala 200:20]
  reg  signs_1_8; // @[block_division.scala 200:20]
  reg  signs_1_9; // @[block_division.scala 200:20]
  reg  signs_1_10; // @[block_division.scala 200:20]
  reg  signs_1_11; // @[block_division.scala 200:20]
  reg  signs_1_12; // @[block_division.scala 200:20]
  reg  signs_1_13; // @[block_division.scala 200:20]
  reg  signs_1_14; // @[block_division.scala 200:20]
  reg  signs_1_15; // @[block_division.scala 200:20]
  reg  signs_1_16; // @[block_division.scala 200:20]
  reg  signs_1_17; // @[block_division.scala 200:20]
  reg  signs_1_18; // @[block_division.scala 200:20]
  reg  signs_1_19; // @[block_division.scala 200:20]
  reg  signs_1_20; // @[block_division.scala 200:20]
  reg  signs_1_21; // @[block_division.scala 200:20]
  reg  signs_1_22; // @[block_division.scala 200:20]
  reg  signs_1_23; // @[block_division.scala 200:20]
  reg  signs_1_24; // @[block_division.scala 200:20]
  reg  signs_1_25; // @[block_division.scala 200:20]
  reg  signs_1_26; // @[block_division.scala 200:20]
  reg  signs_1_27; // @[block_division.scala 200:20]
  reg  signs_1_28; // @[block_division.scala 200:20]
  reg  signs_1_29; // @[block_division.scala 200:20]
  reg  signs_1_30; // @[block_division.scala 200:20]
  reg  signs_1_31; // @[block_division.scala 200:20]
  reg  signs_1_32; // @[block_division.scala 200:20]
  reg  signs_1_33; // @[block_division.scala 200:20]
  reg  signs_1_34; // @[block_division.scala 200:20]
  reg  signs_1_35; // @[block_division.scala 200:20]
  reg  signs_1_36; // @[block_division.scala 200:20]
  reg  signs_1_37; // @[block_division.scala 200:20]
  reg  signs_1_38; // @[block_division.scala 200:20]
  reg  signs_1_39; // @[block_division.scala 200:20]
  reg  signs_1_40; // @[block_division.scala 200:20]
  reg  signs_1_41; // @[block_division.scala 200:20]
  reg  signs_1_42; // @[block_division.scala 200:20]
  reg  signs_1_43; // @[block_division.scala 200:20]
  reg  signs_1_44; // @[block_division.scala 200:20]
  reg  signs_1_45; // @[block_division.scala 200:20]
  reg  signs_1_46; // @[block_division.scala 200:20]
  reg  signs_1_47; // @[block_division.scala 200:20]
  reg  signs_1_48; // @[block_division.scala 200:20]
  reg  signs_1_49; // @[block_division.scala 200:20]
  reg  signs_1_50; // @[block_division.scala 200:20]
  reg  signs_1_51; // @[block_division.scala 200:20]
  reg  signs_1_52; // @[block_division.scala 200:20]
  reg  signs_1_53; // @[block_division.scala 200:20]
  reg  signs_1_54; // @[block_division.scala 200:20]
  reg  signs_1_55; // @[block_division.scala 200:20]
  reg  signs_1_56; // @[block_division.scala 200:20]
  reg  signs_1_57; // @[block_division.scala 200:20]
  reg  signs_1_58; // @[block_division.scala 200:20]
  reg  signs_1_59; // @[block_division.scala 200:20]
  reg  signs_1_60; // @[block_division.scala 200:20]
  reg  signs_1_61; // @[block_division.scala 200:20]
  reg  signs_1_62; // @[block_division.scala 200:20]
  reg  signs_1_63; // @[block_division.scala 200:20]
  reg [5:0] two_complement_1_0; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_1; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_2; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_3; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_4; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_5; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_6; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_7; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_8; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_9; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_10; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_11; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_12; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_13; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_14; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_15; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_16; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_17; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_18; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_19; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_20; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_21; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_22; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_23; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_24; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_25; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_26; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_27; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_28; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_29; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_30; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_31; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_32; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_33; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_34; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_35; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_36; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_37; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_38; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_39; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_40; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_41; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_42; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_43; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_44; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_45; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_46; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_47; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_48; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_49; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_50; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_51; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_52; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_53; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_54; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_55; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_56; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_57; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_58; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_59; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_60; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_61; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_62; // @[block_division.scala 201:29]
  reg [5:0] two_complement_1_63; // @[block_division.scala 201:29]
  reg [5:0] two_complement_buffer_1_0; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_1; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_2; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_3; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_4; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_5; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_6; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_7; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_8; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_9; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_10; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_11; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_12; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_13; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_14; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_15; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_16; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_17; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_18; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_19; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_20; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_21; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_22; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_23; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_24; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_25; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_26; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_27; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_28; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_29; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_30; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_31; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_32; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_33; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_34; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_35; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_36; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_37; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_38; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_39; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_40; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_41; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_42; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_43; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_44; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_45; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_46; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_47; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_48; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_49; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_50; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_51; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_52; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_53; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_54; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_55; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_56; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_57; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_58; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_59; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_60; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_61; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_62; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_1_63; // @[block_division.scala 202:36]
  reg [4:0] multiplierReg_64; // @[block_division.scala 204:34]
  reg  signReg_64; // @[block_division.scala 205:28]
  wire [9:0] multiplication_64 = multiplierReg_64 * io_man_b_64; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_0_T_11 = multiplication_64 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_64; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_0_T_8 = {1'h0,dotProductRegs_1_0}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_0_T_9 = ~_two_complement_0_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_0_T_11 = _two_complement_0_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_65; // @[block_division.scala 204:34]
  reg  signReg_65; // @[block_division.scala 205:28]
  wire [9:0] multiplication_65 = multiplierReg_65 * io_man_b_65; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_1_T_11 = multiplication_65 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_65; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_1_T_8 = {1'h0,dotProductRegs_1_1}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_1_T_9 = ~_two_complement_1_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_1_T_11 = _two_complement_1_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_66; // @[block_division.scala 204:34]
  reg  signReg_66; // @[block_division.scala 205:28]
  wire [9:0] multiplication_66 = multiplierReg_66 * io_man_b_66; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_2_T_11 = multiplication_66 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_66; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_2_T_8 = {1'h0,dotProductRegs_1_2}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_2_T_9 = ~_two_complement_2_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_2_T_11 = _two_complement_2_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_67; // @[block_division.scala 204:34]
  reg  signReg_67; // @[block_division.scala 205:28]
  wire [9:0] multiplication_67 = multiplierReg_67 * io_man_b_67; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_3_T_11 = multiplication_67 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_67; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_3_T_8 = {1'h0,dotProductRegs_1_3}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_3_T_9 = ~_two_complement_3_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_3_T_11 = _two_complement_3_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_68; // @[block_division.scala 204:34]
  reg  signReg_68; // @[block_division.scala 205:28]
  wire [9:0] multiplication_68 = multiplierReg_68 * io_man_b_68; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_4_T_11 = multiplication_68 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_68; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_4_T_8 = {1'h0,dotProductRegs_1_4}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_4_T_9 = ~_two_complement_4_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_4_T_11 = _two_complement_4_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_69; // @[block_division.scala 204:34]
  reg  signReg_69; // @[block_division.scala 205:28]
  wire [9:0] multiplication_69 = multiplierReg_69 * io_man_b_69; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_5_T_11 = multiplication_69 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_69; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_5_T_8 = {1'h0,dotProductRegs_1_5}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_5_T_9 = ~_two_complement_5_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_5_T_11 = _two_complement_5_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_70; // @[block_division.scala 204:34]
  reg  signReg_70; // @[block_division.scala 205:28]
  wire [9:0] multiplication_70 = multiplierReg_70 * io_man_b_70; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_6_T_11 = multiplication_70 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_70; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_6_T_8 = {1'h0,dotProductRegs_1_6}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_6_T_9 = ~_two_complement_6_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_6_T_11 = _two_complement_6_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_71; // @[block_division.scala 204:34]
  reg  signReg_71; // @[block_division.scala 205:28]
  wire [9:0] multiplication_71 = multiplierReg_71 * io_man_b_71; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_7_T_11 = multiplication_71 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_71; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_7_T_8 = {1'h0,dotProductRegs_1_7}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_7_T_9 = ~_two_complement_7_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_7_T_11 = _two_complement_7_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_72; // @[block_division.scala 204:34]
  reg  signReg_72; // @[block_division.scala 205:28]
  wire [9:0] multiplication_72 = multiplierReg_72 * io_man_b_72; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_8_T_11 = multiplication_72 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_72; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_8_T_8 = {1'h0,dotProductRegs_1_8}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_8_T_9 = ~_two_complement_8_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_8_T_11 = _two_complement_8_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_73; // @[block_division.scala 204:34]
  reg  signReg_73; // @[block_division.scala 205:28]
  wire [9:0] multiplication_73 = multiplierReg_73 * io_man_b_73; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_9_T_11 = multiplication_73 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_73; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_9_T_8 = {1'h0,dotProductRegs_1_9}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_9_T_9 = ~_two_complement_9_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_9_T_11 = _two_complement_9_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_74; // @[block_division.scala 204:34]
  reg  signReg_74; // @[block_division.scala 205:28]
  wire [9:0] multiplication_74 = multiplierReg_74 * io_man_b_74; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_10_T_11 = multiplication_74 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_74; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_10_T_8 = {1'h0,dotProductRegs_1_10}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_10_T_9 = ~_two_complement_10_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_10_T_11 = _two_complement_10_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_75; // @[block_division.scala 204:34]
  reg  signReg_75; // @[block_division.scala 205:28]
  wire [9:0] multiplication_75 = multiplierReg_75 * io_man_b_75; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_11_T_11 = multiplication_75 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_75; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_11_T_8 = {1'h0,dotProductRegs_1_11}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_11_T_9 = ~_two_complement_11_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_11_T_11 = _two_complement_11_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_76; // @[block_division.scala 204:34]
  reg  signReg_76; // @[block_division.scala 205:28]
  wire [9:0] multiplication_76 = multiplierReg_76 * io_man_b_76; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_12_T_11 = multiplication_76 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_76; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_12_T_8 = {1'h0,dotProductRegs_1_12}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_12_T_9 = ~_two_complement_12_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_12_T_11 = _two_complement_12_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_77; // @[block_division.scala 204:34]
  reg  signReg_77; // @[block_division.scala 205:28]
  wire [9:0] multiplication_77 = multiplierReg_77 * io_man_b_77; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_13_T_11 = multiplication_77 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_77; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_13_T_8 = {1'h0,dotProductRegs_1_13}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_13_T_9 = ~_two_complement_13_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_13_T_11 = _two_complement_13_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_78; // @[block_division.scala 204:34]
  reg  signReg_78; // @[block_division.scala 205:28]
  wire [9:0] multiplication_78 = multiplierReg_78 * io_man_b_78; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_14_T_11 = multiplication_78 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_78; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_14_T_8 = {1'h0,dotProductRegs_1_14}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_14_T_9 = ~_two_complement_14_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_14_T_11 = _two_complement_14_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_79; // @[block_division.scala 204:34]
  reg  signReg_79; // @[block_division.scala 205:28]
  wire [9:0] multiplication_79 = multiplierReg_79 * io_man_b_79; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_15_T_11 = multiplication_79 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_79; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_15_T_8 = {1'h0,dotProductRegs_1_15}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_15_T_9 = ~_two_complement_15_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_15_T_11 = _two_complement_15_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_80; // @[block_division.scala 204:34]
  reg  signReg_80; // @[block_division.scala 205:28]
  wire [9:0] multiplication_80 = multiplierReg_80 * io_man_b_80; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_16_T_11 = multiplication_80 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_80; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_16_T_8 = {1'h0,dotProductRegs_1_16}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_16_T_9 = ~_two_complement_16_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_16_T_11 = _two_complement_16_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_81; // @[block_division.scala 204:34]
  reg  signReg_81; // @[block_division.scala 205:28]
  wire [9:0] multiplication_81 = multiplierReg_81 * io_man_b_81; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_17_T_11 = multiplication_81 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_81; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_17_T_8 = {1'h0,dotProductRegs_1_17}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_17_T_9 = ~_two_complement_17_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_17_T_11 = _two_complement_17_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_82; // @[block_division.scala 204:34]
  reg  signReg_82; // @[block_division.scala 205:28]
  wire [9:0] multiplication_82 = multiplierReg_82 * io_man_b_82; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_18_T_11 = multiplication_82 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_82; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_18_T_8 = {1'h0,dotProductRegs_1_18}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_18_T_9 = ~_two_complement_18_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_18_T_11 = _two_complement_18_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_83; // @[block_division.scala 204:34]
  reg  signReg_83; // @[block_division.scala 205:28]
  wire [9:0] multiplication_83 = multiplierReg_83 * io_man_b_83; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_19_T_11 = multiplication_83 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_83; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_19_T_8 = {1'h0,dotProductRegs_1_19}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_19_T_9 = ~_two_complement_19_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_19_T_11 = _two_complement_19_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_84; // @[block_division.scala 204:34]
  reg  signReg_84; // @[block_division.scala 205:28]
  wire [9:0] multiplication_84 = multiplierReg_84 * io_man_b_84; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_20_T_11 = multiplication_84 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_84; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_20_T_8 = {1'h0,dotProductRegs_1_20}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_20_T_9 = ~_two_complement_20_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_20_T_11 = _two_complement_20_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_85; // @[block_division.scala 204:34]
  reg  signReg_85; // @[block_division.scala 205:28]
  wire [9:0] multiplication_85 = multiplierReg_85 * io_man_b_85; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_21_T_11 = multiplication_85 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_85; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_21_T_8 = {1'h0,dotProductRegs_1_21}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_21_T_9 = ~_two_complement_21_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_21_T_11 = _two_complement_21_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_86; // @[block_division.scala 204:34]
  reg  signReg_86; // @[block_division.scala 205:28]
  wire [9:0] multiplication_86 = multiplierReg_86 * io_man_b_86; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_22_T_11 = multiplication_86 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_86; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_22_T_8 = {1'h0,dotProductRegs_1_22}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_22_T_9 = ~_two_complement_22_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_22_T_11 = _two_complement_22_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_87; // @[block_division.scala 204:34]
  reg  signReg_87; // @[block_division.scala 205:28]
  wire [9:0] multiplication_87 = multiplierReg_87 * io_man_b_87; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_23_T_11 = multiplication_87 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_87; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_23_T_8 = {1'h0,dotProductRegs_1_23}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_23_T_9 = ~_two_complement_23_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_23_T_11 = _two_complement_23_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_88; // @[block_division.scala 204:34]
  reg  signReg_88; // @[block_division.scala 205:28]
  wire [9:0] multiplication_88 = multiplierReg_88 * io_man_b_88; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_24_T_11 = multiplication_88 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_88; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_24_T_8 = {1'h0,dotProductRegs_1_24}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_24_T_9 = ~_two_complement_24_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_24_T_11 = _two_complement_24_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_89; // @[block_division.scala 204:34]
  reg  signReg_89; // @[block_division.scala 205:28]
  wire [9:0] multiplication_89 = multiplierReg_89 * io_man_b_89; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_25_T_11 = multiplication_89 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_89; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_25_T_8 = {1'h0,dotProductRegs_1_25}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_25_T_9 = ~_two_complement_25_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_25_T_11 = _two_complement_25_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_90; // @[block_division.scala 204:34]
  reg  signReg_90; // @[block_division.scala 205:28]
  wire [9:0] multiplication_90 = multiplierReg_90 * io_man_b_90; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_26_T_11 = multiplication_90 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_90; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_26_T_8 = {1'h0,dotProductRegs_1_26}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_26_T_9 = ~_two_complement_26_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_26_T_11 = _two_complement_26_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_91; // @[block_division.scala 204:34]
  reg  signReg_91; // @[block_division.scala 205:28]
  wire [9:0] multiplication_91 = multiplierReg_91 * io_man_b_91; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_27_T_11 = multiplication_91 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_91; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_27_T_8 = {1'h0,dotProductRegs_1_27}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_27_T_9 = ~_two_complement_27_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_27_T_11 = _two_complement_27_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_92; // @[block_division.scala 204:34]
  reg  signReg_92; // @[block_division.scala 205:28]
  wire [9:0] multiplication_92 = multiplierReg_92 * io_man_b_92; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_28_T_11 = multiplication_92 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_92; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_28_T_8 = {1'h0,dotProductRegs_1_28}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_28_T_9 = ~_two_complement_28_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_28_T_11 = _two_complement_28_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_93; // @[block_division.scala 204:34]
  reg  signReg_93; // @[block_division.scala 205:28]
  wire [9:0] multiplication_93 = multiplierReg_93 * io_man_b_93; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_29_T_11 = multiplication_93 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_93; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_29_T_8 = {1'h0,dotProductRegs_1_29}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_29_T_9 = ~_two_complement_29_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_29_T_11 = _two_complement_29_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_94; // @[block_division.scala 204:34]
  reg  signReg_94; // @[block_division.scala 205:28]
  wire [9:0] multiplication_94 = multiplierReg_94 * io_man_b_94; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_30_T_11 = multiplication_94 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_94; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_30_T_8 = {1'h0,dotProductRegs_1_30}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_30_T_9 = ~_two_complement_30_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_30_T_11 = _two_complement_30_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_95; // @[block_division.scala 204:34]
  reg  signReg_95; // @[block_division.scala 205:28]
  wire [9:0] multiplication_95 = multiplierReg_95 * io_man_b_95; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_31_T_11 = multiplication_95 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_95; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_31_T_8 = {1'h0,dotProductRegs_1_31}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_31_T_9 = ~_two_complement_31_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_31_T_11 = _two_complement_31_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_96; // @[block_division.scala 204:34]
  reg  signReg_96; // @[block_division.scala 205:28]
  wire [9:0] multiplication_96 = multiplierReg_96 * io_man_b_96; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_32_T_11 = multiplication_96 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_96; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_32_T_8 = {1'h0,dotProductRegs_1_32}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_32_T_9 = ~_two_complement_32_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_32_T_11 = _two_complement_32_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_97; // @[block_division.scala 204:34]
  reg  signReg_97; // @[block_division.scala 205:28]
  wire [9:0] multiplication_97 = multiplierReg_97 * io_man_b_97; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_33_T_11 = multiplication_97 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_97; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_33_T_8 = {1'h0,dotProductRegs_1_33}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_33_T_9 = ~_two_complement_33_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_33_T_11 = _two_complement_33_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_98; // @[block_division.scala 204:34]
  reg  signReg_98; // @[block_division.scala 205:28]
  wire [9:0] multiplication_98 = multiplierReg_98 * io_man_b_98; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_34_T_11 = multiplication_98 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_98; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_34_T_8 = {1'h0,dotProductRegs_1_34}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_34_T_9 = ~_two_complement_34_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_34_T_11 = _two_complement_34_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_99; // @[block_division.scala 204:34]
  reg  signReg_99; // @[block_division.scala 205:28]
  wire [9:0] multiplication_99 = multiplierReg_99 * io_man_b_99; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_35_T_11 = multiplication_99 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_99; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_35_T_8 = {1'h0,dotProductRegs_1_35}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_35_T_9 = ~_two_complement_35_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_35_T_11 = _two_complement_35_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_100; // @[block_division.scala 204:34]
  reg  signReg_100; // @[block_division.scala 205:28]
  wire [9:0] multiplication_100 = multiplierReg_100 * io_man_b_100; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_36_T_11 = multiplication_100 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_100; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_36_T_8 = {1'h0,dotProductRegs_1_36}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_36_T_9 = ~_two_complement_36_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_36_T_11 = _two_complement_36_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_101; // @[block_division.scala 204:34]
  reg  signReg_101; // @[block_division.scala 205:28]
  wire [9:0] multiplication_101 = multiplierReg_101 * io_man_b_101; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_37_T_11 = multiplication_101 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_101; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_37_T_8 = {1'h0,dotProductRegs_1_37}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_37_T_9 = ~_two_complement_37_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_37_T_11 = _two_complement_37_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_102; // @[block_division.scala 204:34]
  reg  signReg_102; // @[block_division.scala 205:28]
  wire [9:0] multiplication_102 = multiplierReg_102 * io_man_b_102; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_38_T_11 = multiplication_102 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_102; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_38_T_8 = {1'h0,dotProductRegs_1_38}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_38_T_9 = ~_two_complement_38_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_38_T_11 = _two_complement_38_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_103; // @[block_division.scala 204:34]
  reg  signReg_103; // @[block_division.scala 205:28]
  wire [9:0] multiplication_103 = multiplierReg_103 * io_man_b_103; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_39_T_11 = multiplication_103 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_103; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_39_T_8 = {1'h0,dotProductRegs_1_39}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_39_T_9 = ~_two_complement_39_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_39_T_11 = _two_complement_39_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_104; // @[block_division.scala 204:34]
  reg  signReg_104; // @[block_division.scala 205:28]
  wire [9:0] multiplication_104 = multiplierReg_104 * io_man_b_104; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_40_T_11 = multiplication_104 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_104; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_40_T_8 = {1'h0,dotProductRegs_1_40}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_40_T_9 = ~_two_complement_40_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_40_T_11 = _two_complement_40_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_105; // @[block_division.scala 204:34]
  reg  signReg_105; // @[block_division.scala 205:28]
  wire [9:0] multiplication_105 = multiplierReg_105 * io_man_b_105; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_41_T_11 = multiplication_105 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_105; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_41_T_8 = {1'h0,dotProductRegs_1_41}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_41_T_9 = ~_two_complement_41_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_41_T_11 = _two_complement_41_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_106; // @[block_division.scala 204:34]
  reg  signReg_106; // @[block_division.scala 205:28]
  wire [9:0] multiplication_106 = multiplierReg_106 * io_man_b_106; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_42_T_11 = multiplication_106 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_106; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_42_T_8 = {1'h0,dotProductRegs_1_42}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_42_T_9 = ~_two_complement_42_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_42_T_11 = _two_complement_42_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_107; // @[block_division.scala 204:34]
  reg  signReg_107; // @[block_division.scala 205:28]
  wire [9:0] multiplication_107 = multiplierReg_107 * io_man_b_107; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_43_T_11 = multiplication_107 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_107; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_43_T_8 = {1'h0,dotProductRegs_1_43}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_43_T_9 = ~_two_complement_43_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_43_T_11 = _two_complement_43_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_108; // @[block_division.scala 204:34]
  reg  signReg_108; // @[block_division.scala 205:28]
  wire [9:0] multiplication_108 = multiplierReg_108 * io_man_b_108; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_44_T_11 = multiplication_108 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_108; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_44_T_8 = {1'h0,dotProductRegs_1_44}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_44_T_9 = ~_two_complement_44_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_44_T_11 = _two_complement_44_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_109; // @[block_division.scala 204:34]
  reg  signReg_109; // @[block_division.scala 205:28]
  wire [9:0] multiplication_109 = multiplierReg_109 * io_man_b_109; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_45_T_11 = multiplication_109 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_109; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_45_T_8 = {1'h0,dotProductRegs_1_45}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_45_T_9 = ~_two_complement_45_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_45_T_11 = _two_complement_45_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_110; // @[block_division.scala 204:34]
  reg  signReg_110; // @[block_division.scala 205:28]
  wire [9:0] multiplication_110 = multiplierReg_110 * io_man_b_110; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_46_T_11 = multiplication_110 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_110; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_46_T_8 = {1'h0,dotProductRegs_1_46}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_46_T_9 = ~_two_complement_46_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_46_T_11 = _two_complement_46_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_111; // @[block_division.scala 204:34]
  reg  signReg_111; // @[block_division.scala 205:28]
  wire [9:0] multiplication_111 = multiplierReg_111 * io_man_b_111; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_47_T_11 = multiplication_111 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_111; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_47_T_8 = {1'h0,dotProductRegs_1_47}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_47_T_9 = ~_two_complement_47_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_47_T_11 = _two_complement_47_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_112; // @[block_division.scala 204:34]
  reg  signReg_112; // @[block_division.scala 205:28]
  wire [9:0] multiplication_112 = multiplierReg_112 * io_man_b_112; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_48_T_11 = multiplication_112 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_112; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_48_T_8 = {1'h0,dotProductRegs_1_48}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_48_T_9 = ~_two_complement_48_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_48_T_11 = _two_complement_48_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_113; // @[block_division.scala 204:34]
  reg  signReg_113; // @[block_division.scala 205:28]
  wire [9:0] multiplication_113 = multiplierReg_113 * io_man_b_113; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_49_T_11 = multiplication_113 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_113; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_49_T_8 = {1'h0,dotProductRegs_1_49}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_49_T_9 = ~_two_complement_49_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_49_T_11 = _two_complement_49_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_114; // @[block_division.scala 204:34]
  reg  signReg_114; // @[block_division.scala 205:28]
  wire [9:0] multiplication_114 = multiplierReg_114 * io_man_b_114; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_50_T_11 = multiplication_114 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_114; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_50_T_8 = {1'h0,dotProductRegs_1_50}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_50_T_9 = ~_two_complement_50_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_50_T_11 = _two_complement_50_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_115; // @[block_division.scala 204:34]
  reg  signReg_115; // @[block_division.scala 205:28]
  wire [9:0] multiplication_115 = multiplierReg_115 * io_man_b_115; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_51_T_11 = multiplication_115 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_115; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_51_T_8 = {1'h0,dotProductRegs_1_51}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_51_T_9 = ~_two_complement_51_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_51_T_11 = _two_complement_51_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_116; // @[block_division.scala 204:34]
  reg  signReg_116; // @[block_division.scala 205:28]
  wire [9:0] multiplication_116 = multiplierReg_116 * io_man_b_116; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_52_T_11 = multiplication_116 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_116; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_52_T_8 = {1'h0,dotProductRegs_1_52}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_52_T_9 = ~_two_complement_52_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_52_T_11 = _two_complement_52_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_117; // @[block_division.scala 204:34]
  reg  signReg_117; // @[block_division.scala 205:28]
  wire [9:0] multiplication_117 = multiplierReg_117 * io_man_b_117; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_53_T_11 = multiplication_117 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_117; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_53_T_8 = {1'h0,dotProductRegs_1_53}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_53_T_9 = ~_two_complement_53_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_53_T_11 = _two_complement_53_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_118; // @[block_division.scala 204:34]
  reg  signReg_118; // @[block_division.scala 205:28]
  wire [9:0] multiplication_118 = multiplierReg_118 * io_man_b_118; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_54_T_11 = multiplication_118 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_118; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_54_T_8 = {1'h0,dotProductRegs_1_54}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_54_T_9 = ~_two_complement_54_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_54_T_11 = _two_complement_54_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_119; // @[block_division.scala 204:34]
  reg  signReg_119; // @[block_division.scala 205:28]
  wire [9:0] multiplication_119 = multiplierReg_119 * io_man_b_119; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_55_T_11 = multiplication_119 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_119; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_55_T_8 = {1'h0,dotProductRegs_1_55}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_55_T_9 = ~_two_complement_55_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_55_T_11 = _two_complement_55_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_120; // @[block_division.scala 204:34]
  reg  signReg_120; // @[block_division.scala 205:28]
  wire [9:0] multiplication_120 = multiplierReg_120 * io_man_b_120; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_56_T_11 = multiplication_120 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_120; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_56_T_8 = {1'h0,dotProductRegs_1_56}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_56_T_9 = ~_two_complement_56_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_56_T_11 = _two_complement_56_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_121; // @[block_division.scala 204:34]
  reg  signReg_121; // @[block_division.scala 205:28]
  wire [9:0] multiplication_121 = multiplierReg_121 * io_man_b_121; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_57_T_11 = multiplication_121 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_121; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_57_T_8 = {1'h0,dotProductRegs_1_57}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_57_T_9 = ~_two_complement_57_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_57_T_11 = _two_complement_57_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_122; // @[block_division.scala 204:34]
  reg  signReg_122; // @[block_division.scala 205:28]
  wire [9:0] multiplication_122 = multiplierReg_122 * io_man_b_122; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_58_T_11 = multiplication_122 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_122; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_58_T_8 = {1'h0,dotProductRegs_1_58}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_58_T_9 = ~_two_complement_58_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_58_T_11 = _two_complement_58_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_123; // @[block_division.scala 204:34]
  reg  signReg_123; // @[block_division.scala 205:28]
  wire [9:0] multiplication_123 = multiplierReg_123 * io_man_b_123; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_59_T_11 = multiplication_123 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_123; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_59_T_8 = {1'h0,dotProductRegs_1_59}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_59_T_9 = ~_two_complement_59_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_59_T_11 = _two_complement_59_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_124; // @[block_division.scala 204:34]
  reg  signReg_124; // @[block_division.scala 205:28]
  wire [9:0] multiplication_124 = multiplierReg_124 * io_man_b_124; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_60_T_11 = multiplication_124 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_124; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_60_T_8 = {1'h0,dotProductRegs_1_60}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_60_T_9 = ~_two_complement_60_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_60_T_11 = _two_complement_60_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_125; // @[block_division.scala 204:34]
  reg  signReg_125; // @[block_division.scala 205:28]
  wire [9:0] multiplication_125 = multiplierReg_125 * io_man_b_125; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_61_T_11 = multiplication_125 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_125; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_61_T_8 = {1'h0,dotProductRegs_1_61}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_61_T_9 = ~_two_complement_61_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_61_T_11 = _two_complement_61_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_126; // @[block_division.scala 204:34]
  reg  signReg_126; // @[block_division.scala 205:28]
  wire [9:0] multiplication_126 = multiplierReg_126 * io_man_b_126; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_62_T_11 = multiplication_126 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_126; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_62_T_8 = {1'h0,dotProductRegs_1_62}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_62_T_9 = ~_two_complement_62_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_62_T_11 = _two_complement_62_T_9 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_127; // @[block_division.scala 204:34]
  reg  signReg_127; // @[block_division.scala 205:28]
  wire [9:0] multiplication_127 = multiplierReg_127 * io_man_b_127; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_63_T_11 = multiplication_127 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_127; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_63_T_8 = {1'h0,dotProductRegs_1_63}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_63_T_9 = ~_two_complement_63_T_8; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_63_T_11 = _two_complement_63_T_9 + 6'h1; // @[block_division.scala 213:38]
  wire [6:0] _sum_T_62 = $signed(two_complement_buffer_1_0) + $signed(two_complement_buffer_1_1); // @[block_division.scala 218:46]
  wire [6:0] _GEN_192 = {{1{two_complement_buffer_1_2[5]}},two_complement_buffer_1_2}; // @[block_division.scala 218:46]
  wire [7:0] _sum_T_63 = $signed(_sum_T_62) + $signed(_GEN_192); // @[block_division.scala 218:46]
  wire [7:0] _GEN_193 = {{2{two_complement_buffer_1_3[5]}},two_complement_buffer_1_3}; // @[block_division.scala 218:46]
  wire [8:0] _sum_T_64 = $signed(_sum_T_63) + $signed(_GEN_193); // @[block_division.scala 218:46]
  wire [8:0] _GEN_194 = {{3{two_complement_buffer_1_4[5]}},two_complement_buffer_1_4}; // @[block_division.scala 218:46]
  wire [9:0] _sum_T_65 = $signed(_sum_T_64) + $signed(_GEN_194); // @[block_division.scala 218:46]
  wire [9:0] _GEN_195 = {{4{two_complement_buffer_1_5[5]}},two_complement_buffer_1_5}; // @[block_division.scala 218:46]
  wire [10:0] _sum_T_66 = $signed(_sum_T_65) + $signed(_GEN_195); // @[block_division.scala 218:46]
  wire [10:0] _GEN_196 = {{5{two_complement_buffer_1_6[5]}},two_complement_buffer_1_6}; // @[block_division.scala 218:46]
  wire [11:0] _sum_T_67 = $signed(_sum_T_66) + $signed(_GEN_196); // @[block_division.scala 218:46]
  wire [11:0] _GEN_197 = {{6{two_complement_buffer_1_7[5]}},two_complement_buffer_1_7}; // @[block_division.scala 218:46]
  wire [12:0] _sum_T_68 = $signed(_sum_T_67) + $signed(_GEN_197); // @[block_division.scala 218:46]
  wire [12:0] _GEN_198 = {{7{two_complement_buffer_1_8[5]}},two_complement_buffer_1_8}; // @[block_division.scala 218:46]
  wire [13:0] _sum_T_69 = $signed(_sum_T_68) + $signed(_GEN_198); // @[block_division.scala 218:46]
  wire [13:0] _GEN_199 = {{8{two_complement_buffer_1_9[5]}},two_complement_buffer_1_9}; // @[block_division.scala 218:46]
  wire [14:0] _sum_T_70 = $signed(_sum_T_69) + $signed(_GEN_199); // @[block_division.scala 218:46]
  wire [14:0] _GEN_200 = {{9{two_complement_buffer_1_10[5]}},two_complement_buffer_1_10}; // @[block_division.scala 218:46]
  wire [15:0] _sum_T_71 = $signed(_sum_T_70) + $signed(_GEN_200); // @[block_division.scala 218:46]
  wire [15:0] _GEN_201 = {{10{two_complement_buffer_1_11[5]}},two_complement_buffer_1_11}; // @[block_division.scala 218:46]
  wire [16:0] _sum_T_72 = $signed(_sum_T_71) + $signed(_GEN_201); // @[block_division.scala 218:46]
  wire [16:0] _GEN_202 = {{11{two_complement_buffer_1_12[5]}},two_complement_buffer_1_12}; // @[block_division.scala 218:46]
  wire [17:0] _sum_T_73 = $signed(_sum_T_72) + $signed(_GEN_202); // @[block_division.scala 218:46]
  wire [17:0] _GEN_203 = {{12{two_complement_buffer_1_13[5]}},two_complement_buffer_1_13}; // @[block_division.scala 218:46]
  wire [18:0] _sum_T_74 = $signed(_sum_T_73) + $signed(_GEN_203); // @[block_division.scala 218:46]
  wire [18:0] _GEN_204 = {{13{two_complement_buffer_1_14[5]}},two_complement_buffer_1_14}; // @[block_division.scala 218:46]
  wire [19:0] _sum_T_75 = $signed(_sum_T_74) + $signed(_GEN_204); // @[block_division.scala 218:46]
  wire [19:0] _GEN_205 = {{14{two_complement_buffer_1_15[5]}},two_complement_buffer_1_15}; // @[block_division.scala 218:46]
  wire [20:0] _sum_T_76 = $signed(_sum_T_75) + $signed(_GEN_205); // @[block_division.scala 218:46]
  wire [20:0] _GEN_206 = {{15{two_complement_buffer_1_16[5]}},two_complement_buffer_1_16}; // @[block_division.scala 218:46]
  wire [21:0] _sum_T_77 = $signed(_sum_T_76) + $signed(_GEN_206); // @[block_division.scala 218:46]
  wire [21:0] _GEN_207 = {{16{two_complement_buffer_1_17[5]}},two_complement_buffer_1_17}; // @[block_division.scala 218:46]
  wire [22:0] _sum_T_78 = $signed(_sum_T_77) + $signed(_GEN_207); // @[block_division.scala 218:46]
  wire [22:0] _GEN_208 = {{17{two_complement_buffer_1_18[5]}},two_complement_buffer_1_18}; // @[block_division.scala 218:46]
  wire [23:0] _sum_T_79 = $signed(_sum_T_78) + $signed(_GEN_208); // @[block_division.scala 218:46]
  wire [23:0] _GEN_209 = {{18{two_complement_buffer_1_19[5]}},two_complement_buffer_1_19}; // @[block_division.scala 218:46]
  wire [24:0] _sum_T_80 = $signed(_sum_T_79) + $signed(_GEN_209); // @[block_division.scala 218:46]
  wire [24:0] _GEN_210 = {{19{two_complement_buffer_1_20[5]}},two_complement_buffer_1_20}; // @[block_division.scala 218:46]
  wire [25:0] _sum_T_81 = $signed(_sum_T_80) + $signed(_GEN_210); // @[block_division.scala 218:46]
  wire [25:0] _GEN_211 = {{20{two_complement_buffer_1_21[5]}},two_complement_buffer_1_21}; // @[block_division.scala 218:46]
  wire [26:0] _sum_T_82 = $signed(_sum_T_81) + $signed(_GEN_211); // @[block_division.scala 218:46]
  wire [26:0] _GEN_212 = {{21{two_complement_buffer_1_22[5]}},two_complement_buffer_1_22}; // @[block_division.scala 218:46]
  wire [27:0] _sum_T_83 = $signed(_sum_T_82) + $signed(_GEN_212); // @[block_division.scala 218:46]
  wire [27:0] _GEN_213 = {{22{two_complement_buffer_1_23[5]}},two_complement_buffer_1_23}; // @[block_division.scala 218:46]
  wire [28:0] _sum_T_84 = $signed(_sum_T_83) + $signed(_GEN_213); // @[block_division.scala 218:46]
  wire [28:0] _GEN_214 = {{23{two_complement_buffer_1_24[5]}},two_complement_buffer_1_24}; // @[block_division.scala 218:46]
  wire [29:0] _sum_T_85 = $signed(_sum_T_84) + $signed(_GEN_214); // @[block_division.scala 218:46]
  wire [29:0] _GEN_215 = {{24{two_complement_buffer_1_25[5]}},two_complement_buffer_1_25}; // @[block_division.scala 218:46]
  wire [30:0] _sum_T_86 = $signed(_sum_T_85) + $signed(_GEN_215); // @[block_division.scala 218:46]
  wire [30:0] _GEN_216 = {{25{two_complement_buffer_1_26[5]}},two_complement_buffer_1_26}; // @[block_division.scala 218:46]
  wire [31:0] _sum_T_87 = $signed(_sum_T_86) + $signed(_GEN_216); // @[block_division.scala 218:46]
  wire [31:0] _GEN_217 = {{26{two_complement_buffer_1_27[5]}},two_complement_buffer_1_27}; // @[block_division.scala 218:46]
  wire [32:0] _sum_T_88 = $signed(_sum_T_87) + $signed(_GEN_217); // @[block_division.scala 218:46]
  wire [32:0] _GEN_218 = {{27{two_complement_buffer_1_28[5]}},two_complement_buffer_1_28}; // @[block_division.scala 218:46]
  wire [33:0] _sum_T_89 = $signed(_sum_T_88) + $signed(_GEN_218); // @[block_division.scala 218:46]
  wire [33:0] _GEN_219 = {{28{two_complement_buffer_1_29[5]}},two_complement_buffer_1_29}; // @[block_division.scala 218:46]
  wire [34:0] _sum_T_90 = $signed(_sum_T_89) + $signed(_GEN_219); // @[block_division.scala 218:46]
  wire [34:0] _GEN_220 = {{29{two_complement_buffer_1_30[5]}},two_complement_buffer_1_30}; // @[block_division.scala 218:46]
  wire [35:0] _sum_T_91 = $signed(_sum_T_90) + $signed(_GEN_220); // @[block_division.scala 218:46]
  wire [35:0] _GEN_221 = {{30{two_complement_buffer_1_31[5]}},two_complement_buffer_1_31}; // @[block_division.scala 218:46]
  wire [36:0] _sum_T_92 = $signed(_sum_T_91) + $signed(_GEN_221); // @[block_division.scala 218:46]
  wire [36:0] _GEN_222 = {{31{two_complement_buffer_1_32[5]}},two_complement_buffer_1_32}; // @[block_division.scala 218:46]
  wire [37:0] _sum_T_93 = $signed(_sum_T_92) + $signed(_GEN_222); // @[block_division.scala 218:46]
  wire [37:0] _GEN_223 = {{32{two_complement_buffer_1_33[5]}},two_complement_buffer_1_33}; // @[block_division.scala 218:46]
  wire [38:0] _sum_T_94 = $signed(_sum_T_93) + $signed(_GEN_223); // @[block_division.scala 218:46]
  wire [38:0] _GEN_224 = {{33{two_complement_buffer_1_34[5]}},two_complement_buffer_1_34}; // @[block_division.scala 218:46]
  wire [39:0] _sum_T_95 = $signed(_sum_T_94) + $signed(_GEN_224); // @[block_division.scala 218:46]
  wire [39:0] _GEN_225 = {{34{two_complement_buffer_1_35[5]}},two_complement_buffer_1_35}; // @[block_division.scala 218:46]
  wire [40:0] _sum_T_96 = $signed(_sum_T_95) + $signed(_GEN_225); // @[block_division.scala 218:46]
  wire [40:0] _GEN_226 = {{35{two_complement_buffer_1_36[5]}},two_complement_buffer_1_36}; // @[block_division.scala 218:46]
  wire [41:0] _sum_T_97 = $signed(_sum_T_96) + $signed(_GEN_226); // @[block_division.scala 218:46]
  wire [41:0] _GEN_227 = {{36{two_complement_buffer_1_37[5]}},two_complement_buffer_1_37}; // @[block_division.scala 218:46]
  wire [42:0] _sum_T_98 = $signed(_sum_T_97) + $signed(_GEN_227); // @[block_division.scala 218:46]
  wire [42:0] _GEN_228 = {{37{two_complement_buffer_1_38[5]}},two_complement_buffer_1_38}; // @[block_division.scala 218:46]
  wire [43:0] _sum_T_99 = $signed(_sum_T_98) + $signed(_GEN_228); // @[block_division.scala 218:46]
  wire [43:0] _GEN_229 = {{38{two_complement_buffer_1_39[5]}},two_complement_buffer_1_39}; // @[block_division.scala 218:46]
  wire [44:0] _sum_T_100 = $signed(_sum_T_99) + $signed(_GEN_229); // @[block_division.scala 218:46]
  wire [44:0] _GEN_230 = {{39{two_complement_buffer_1_40[5]}},two_complement_buffer_1_40}; // @[block_division.scala 218:46]
  wire [45:0] _sum_T_101 = $signed(_sum_T_100) + $signed(_GEN_230); // @[block_division.scala 218:46]
  wire [45:0] _GEN_231 = {{40{two_complement_buffer_1_41[5]}},two_complement_buffer_1_41}; // @[block_division.scala 218:46]
  wire [46:0] _sum_T_102 = $signed(_sum_T_101) + $signed(_GEN_231); // @[block_division.scala 218:46]
  wire [46:0] _GEN_232 = {{41{two_complement_buffer_1_42[5]}},two_complement_buffer_1_42}; // @[block_division.scala 218:46]
  wire [47:0] _sum_T_103 = $signed(_sum_T_102) + $signed(_GEN_232); // @[block_division.scala 218:46]
  wire [47:0] _GEN_233 = {{42{two_complement_buffer_1_43[5]}},two_complement_buffer_1_43}; // @[block_division.scala 218:46]
  wire [48:0] _sum_T_104 = $signed(_sum_T_103) + $signed(_GEN_233); // @[block_division.scala 218:46]
  wire [48:0] _GEN_234 = {{43{two_complement_buffer_1_44[5]}},two_complement_buffer_1_44}; // @[block_division.scala 218:46]
  wire [49:0] _sum_T_105 = $signed(_sum_T_104) + $signed(_GEN_234); // @[block_division.scala 218:46]
  wire [49:0] _GEN_235 = {{44{two_complement_buffer_1_45[5]}},two_complement_buffer_1_45}; // @[block_division.scala 218:46]
  wire [50:0] _sum_T_106 = $signed(_sum_T_105) + $signed(_GEN_235); // @[block_division.scala 218:46]
  wire [50:0] _GEN_236 = {{45{two_complement_buffer_1_46[5]}},two_complement_buffer_1_46}; // @[block_division.scala 218:46]
  wire [51:0] _sum_T_107 = $signed(_sum_T_106) + $signed(_GEN_236); // @[block_division.scala 218:46]
  wire [51:0] _GEN_237 = {{46{two_complement_buffer_1_47[5]}},two_complement_buffer_1_47}; // @[block_division.scala 218:46]
  wire [52:0] _sum_T_108 = $signed(_sum_T_107) + $signed(_GEN_237); // @[block_division.scala 218:46]
  wire [52:0] _GEN_238 = {{47{two_complement_buffer_1_48[5]}},two_complement_buffer_1_48}; // @[block_division.scala 218:46]
  wire [53:0] _sum_T_109 = $signed(_sum_T_108) + $signed(_GEN_238); // @[block_division.scala 218:46]
  wire [53:0] _GEN_239 = {{48{two_complement_buffer_1_49[5]}},two_complement_buffer_1_49}; // @[block_division.scala 218:46]
  wire [54:0] _sum_T_110 = $signed(_sum_T_109) + $signed(_GEN_239); // @[block_division.scala 218:46]
  wire [54:0] _GEN_240 = {{49{two_complement_buffer_1_50[5]}},two_complement_buffer_1_50}; // @[block_division.scala 218:46]
  wire [55:0] _sum_T_111 = $signed(_sum_T_110) + $signed(_GEN_240); // @[block_division.scala 218:46]
  wire [55:0] _GEN_241 = {{50{two_complement_buffer_1_51[5]}},two_complement_buffer_1_51}; // @[block_division.scala 218:46]
  wire [56:0] _sum_T_112 = $signed(_sum_T_111) + $signed(_GEN_241); // @[block_division.scala 218:46]
  wire [56:0] _GEN_242 = {{51{two_complement_buffer_1_52[5]}},two_complement_buffer_1_52}; // @[block_division.scala 218:46]
  wire [57:0] _sum_T_113 = $signed(_sum_T_112) + $signed(_GEN_242); // @[block_division.scala 218:46]
  wire [57:0] _GEN_243 = {{52{two_complement_buffer_1_53[5]}},two_complement_buffer_1_53}; // @[block_division.scala 218:46]
  wire [58:0] _sum_T_114 = $signed(_sum_T_113) + $signed(_GEN_243); // @[block_division.scala 218:46]
  wire [58:0] _GEN_244 = {{53{two_complement_buffer_1_54[5]}},two_complement_buffer_1_54}; // @[block_division.scala 218:46]
  wire [59:0] _sum_T_115 = $signed(_sum_T_114) + $signed(_GEN_244); // @[block_division.scala 218:46]
  wire [59:0] _GEN_245 = {{54{two_complement_buffer_1_55[5]}},two_complement_buffer_1_55}; // @[block_division.scala 218:46]
  wire [60:0] _sum_T_116 = $signed(_sum_T_115) + $signed(_GEN_245); // @[block_division.scala 218:46]
  wire [60:0] _GEN_246 = {{55{two_complement_buffer_1_56[5]}},two_complement_buffer_1_56}; // @[block_division.scala 218:46]
  wire [61:0] _sum_T_117 = $signed(_sum_T_116) + $signed(_GEN_246); // @[block_division.scala 218:46]
  wire [61:0] _GEN_247 = {{56{two_complement_buffer_1_57[5]}},two_complement_buffer_1_57}; // @[block_division.scala 218:46]
  wire [62:0] _sum_T_118 = $signed(_sum_T_117) + $signed(_GEN_247); // @[block_division.scala 218:46]
  wire [62:0] _GEN_248 = {{57{two_complement_buffer_1_58[5]}},two_complement_buffer_1_58}; // @[block_division.scala 218:46]
  wire [63:0] _sum_T_119 = $signed(_sum_T_118) + $signed(_GEN_248); // @[block_division.scala 218:46]
  wire [63:0] _GEN_249 = {{58{two_complement_buffer_1_59[5]}},two_complement_buffer_1_59}; // @[block_division.scala 218:46]
  wire [64:0] _sum_T_120 = $signed(_sum_T_119) + $signed(_GEN_249); // @[block_division.scala 218:46]
  wire [64:0] _GEN_250 = {{59{two_complement_buffer_1_60[5]}},two_complement_buffer_1_60}; // @[block_division.scala 218:46]
  wire [65:0] _sum_T_121 = $signed(_sum_T_120) + $signed(_GEN_250); // @[block_division.scala 218:46]
  wire [65:0] _GEN_251 = {{60{two_complement_buffer_1_61[5]}},two_complement_buffer_1_61}; // @[block_division.scala 218:46]
  wire [66:0] _sum_T_122 = $signed(_sum_T_121) + $signed(_GEN_251); // @[block_division.scala 218:46]
  wire [66:0] _GEN_252 = {{61{two_complement_buffer_1_62[5]}},two_complement_buffer_1_62}; // @[block_division.scala 218:46]
  wire [67:0] _sum_T_123 = $signed(_sum_T_122) + $signed(_GEN_252); // @[block_division.scala 218:46]
  wire [67:0] _GEN_253 = {{62{two_complement_buffer_1_63[5]}},two_complement_buffer_1_63}; // @[block_division.scala 218:46]
  wire [68:0] sum_1 = $signed(_sum_T_123) + $signed(_GEN_253); // @[block_division.scala 218:46]
  wire [67:0] _acc_1_T_3 = ~sum_1[67:0]; // @[block_division.scala 219:57]
  wire [67:0] _acc_1_T_5 = _acc_1_T_3 + 68'h1; // @[block_division.scala 219:86]
  wire [68:0] _acc_1_T_14 = $signed(_sum_T_123) + $signed(_GEN_253); // @[block_division.scala 219:145]
  wire [68:0] _acc_1_T_15 = _acc_1_T_5 > _GEN_126 ? {{63'd0}, _acc_0_T_13} : _acc_1_T_14; // @[block_division.scala 219:55]
  wire [68:0] _acc_1_T_23 = sum_1[67:0] > _GEN_126 ? {{63'd0}, _dotProductRegs_0_T_1} : _acc_1_T_14; // @[block_division.scala 220:6]
  wire [68:0] _acc_1_T_24 = sum_1[68] ? _acc_1_T_15 : _acc_1_T_23; // @[block_division.scala 219:18]
  wire [8:0] _exp_output_2_T = io_exp_a_2 + io_exp_b_2; // @[block_division.scala 198:34]
  reg [4:0] dotProductRegs_2_0; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_1; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_2; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_3; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_4; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_5; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_6; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_7; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_8; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_9; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_10; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_11; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_12; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_13; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_14; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_15; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_16; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_17; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_18; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_19; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_20; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_21; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_22; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_23; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_24; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_25; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_26; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_27; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_28; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_29; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_30; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_31; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_32; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_33; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_34; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_35; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_36; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_37; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_38; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_39; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_40; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_41; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_42; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_43; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_44; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_45; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_46; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_47; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_48; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_49; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_50; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_51; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_52; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_53; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_54; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_55; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_56; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_57; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_58; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_59; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_60; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_61; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_62; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_2_63; // @[block_division.scala 199:29]
  reg  signs_2_0; // @[block_division.scala 200:20]
  reg  signs_2_1; // @[block_division.scala 200:20]
  reg  signs_2_2; // @[block_division.scala 200:20]
  reg  signs_2_3; // @[block_division.scala 200:20]
  reg  signs_2_4; // @[block_division.scala 200:20]
  reg  signs_2_5; // @[block_division.scala 200:20]
  reg  signs_2_6; // @[block_division.scala 200:20]
  reg  signs_2_7; // @[block_division.scala 200:20]
  reg  signs_2_8; // @[block_division.scala 200:20]
  reg  signs_2_9; // @[block_division.scala 200:20]
  reg  signs_2_10; // @[block_division.scala 200:20]
  reg  signs_2_11; // @[block_division.scala 200:20]
  reg  signs_2_12; // @[block_division.scala 200:20]
  reg  signs_2_13; // @[block_division.scala 200:20]
  reg  signs_2_14; // @[block_division.scala 200:20]
  reg  signs_2_15; // @[block_division.scala 200:20]
  reg  signs_2_16; // @[block_division.scala 200:20]
  reg  signs_2_17; // @[block_division.scala 200:20]
  reg  signs_2_18; // @[block_division.scala 200:20]
  reg  signs_2_19; // @[block_division.scala 200:20]
  reg  signs_2_20; // @[block_division.scala 200:20]
  reg  signs_2_21; // @[block_division.scala 200:20]
  reg  signs_2_22; // @[block_division.scala 200:20]
  reg  signs_2_23; // @[block_division.scala 200:20]
  reg  signs_2_24; // @[block_division.scala 200:20]
  reg  signs_2_25; // @[block_division.scala 200:20]
  reg  signs_2_26; // @[block_division.scala 200:20]
  reg  signs_2_27; // @[block_division.scala 200:20]
  reg  signs_2_28; // @[block_division.scala 200:20]
  reg  signs_2_29; // @[block_division.scala 200:20]
  reg  signs_2_30; // @[block_division.scala 200:20]
  reg  signs_2_31; // @[block_division.scala 200:20]
  reg  signs_2_32; // @[block_division.scala 200:20]
  reg  signs_2_33; // @[block_division.scala 200:20]
  reg  signs_2_34; // @[block_division.scala 200:20]
  reg  signs_2_35; // @[block_division.scala 200:20]
  reg  signs_2_36; // @[block_division.scala 200:20]
  reg  signs_2_37; // @[block_division.scala 200:20]
  reg  signs_2_38; // @[block_division.scala 200:20]
  reg  signs_2_39; // @[block_division.scala 200:20]
  reg  signs_2_40; // @[block_division.scala 200:20]
  reg  signs_2_41; // @[block_division.scala 200:20]
  reg  signs_2_42; // @[block_division.scala 200:20]
  reg  signs_2_43; // @[block_division.scala 200:20]
  reg  signs_2_44; // @[block_division.scala 200:20]
  reg  signs_2_45; // @[block_division.scala 200:20]
  reg  signs_2_46; // @[block_division.scala 200:20]
  reg  signs_2_47; // @[block_division.scala 200:20]
  reg  signs_2_48; // @[block_division.scala 200:20]
  reg  signs_2_49; // @[block_division.scala 200:20]
  reg  signs_2_50; // @[block_division.scala 200:20]
  reg  signs_2_51; // @[block_division.scala 200:20]
  reg  signs_2_52; // @[block_division.scala 200:20]
  reg  signs_2_53; // @[block_division.scala 200:20]
  reg  signs_2_54; // @[block_division.scala 200:20]
  reg  signs_2_55; // @[block_division.scala 200:20]
  reg  signs_2_56; // @[block_division.scala 200:20]
  reg  signs_2_57; // @[block_division.scala 200:20]
  reg  signs_2_58; // @[block_division.scala 200:20]
  reg  signs_2_59; // @[block_division.scala 200:20]
  reg  signs_2_60; // @[block_division.scala 200:20]
  reg  signs_2_61; // @[block_division.scala 200:20]
  reg  signs_2_62; // @[block_division.scala 200:20]
  reg  signs_2_63; // @[block_division.scala 200:20]
  reg [5:0] two_complement_2_0; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_1; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_2; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_3; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_4; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_5; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_6; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_7; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_8; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_9; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_10; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_11; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_12; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_13; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_14; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_15; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_16; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_17; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_18; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_19; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_20; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_21; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_22; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_23; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_24; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_25; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_26; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_27; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_28; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_29; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_30; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_31; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_32; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_33; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_34; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_35; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_36; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_37; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_38; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_39; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_40; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_41; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_42; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_43; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_44; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_45; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_46; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_47; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_48; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_49; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_50; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_51; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_52; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_53; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_54; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_55; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_56; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_57; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_58; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_59; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_60; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_61; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_62; // @[block_division.scala 201:29]
  reg [5:0] two_complement_2_63; // @[block_division.scala 201:29]
  reg [5:0] two_complement_buffer_2_0; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_1; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_2; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_3; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_4; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_5; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_6; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_7; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_8; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_9; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_10; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_11; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_12; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_13; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_14; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_15; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_16; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_17; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_18; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_19; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_20; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_21; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_22; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_23; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_24; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_25; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_26; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_27; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_28; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_29; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_30; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_31; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_32; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_33; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_34; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_35; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_36; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_37; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_38; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_39; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_40; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_41; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_42; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_43; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_44; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_45; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_46; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_47; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_48; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_49; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_50; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_51; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_52; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_53; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_54; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_55; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_56; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_57; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_58; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_59; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_60; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_61; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_62; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_2_63; // @[block_division.scala 202:36]
  reg [4:0] multiplierReg_128; // @[block_division.scala 204:34]
  reg  signReg_128; // @[block_division.scala 205:28]
  wire [9:0] multiplication_128 = multiplierReg_128 * io_man_b_128; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_0_T_17 = multiplication_128 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_128
    ; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_0_T_15 = {1'h0,dotProductRegs_2_0}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_0_T_16 = ~_two_complement_0_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_0_T_18 = _two_complement_0_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_129; // @[block_division.scala 204:34]
  reg  signReg_129; // @[block_division.scala 205:28]
  wire [9:0] multiplication_129 = multiplierReg_129 * io_man_b_129; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_1_T_17 = multiplication_129 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_129
    ; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_1_T_15 = {1'h0,dotProductRegs_2_1}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_1_T_16 = ~_two_complement_1_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_1_T_18 = _two_complement_1_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_130; // @[block_division.scala 204:34]
  reg  signReg_130; // @[block_division.scala 205:28]
  wire [9:0] multiplication_130 = multiplierReg_130 * io_man_b_130; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_2_T_17 = multiplication_130 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_130
    ; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_2_T_15 = {1'h0,dotProductRegs_2_2}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_2_T_16 = ~_two_complement_2_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_2_T_18 = _two_complement_2_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_131; // @[block_division.scala 204:34]
  reg  signReg_131; // @[block_division.scala 205:28]
  wire [9:0] multiplication_131 = multiplierReg_131 * io_man_b_131; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_3_T_17 = multiplication_131 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_131
    ; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_3_T_15 = {1'h0,dotProductRegs_2_3}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_3_T_16 = ~_two_complement_3_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_3_T_18 = _two_complement_3_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_132; // @[block_division.scala 204:34]
  reg  signReg_132; // @[block_division.scala 205:28]
  wire [9:0] multiplication_132 = multiplierReg_132 * io_man_b_132; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_4_T_17 = multiplication_132 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_132
    ; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_4_T_15 = {1'h0,dotProductRegs_2_4}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_4_T_16 = ~_two_complement_4_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_4_T_18 = _two_complement_4_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_133; // @[block_division.scala 204:34]
  reg  signReg_133; // @[block_division.scala 205:28]
  wire [9:0] multiplication_133 = multiplierReg_133 * io_man_b_133; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_5_T_17 = multiplication_133 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_133
    ; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_5_T_15 = {1'h0,dotProductRegs_2_5}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_5_T_16 = ~_two_complement_5_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_5_T_18 = _two_complement_5_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_134; // @[block_division.scala 204:34]
  reg  signReg_134; // @[block_division.scala 205:28]
  wire [9:0] multiplication_134 = multiplierReg_134 * io_man_b_134; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_6_T_17 = multiplication_134 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_134
    ; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_6_T_15 = {1'h0,dotProductRegs_2_6}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_6_T_16 = ~_two_complement_6_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_6_T_18 = _two_complement_6_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_135; // @[block_division.scala 204:34]
  reg  signReg_135; // @[block_division.scala 205:28]
  wire [9:0] multiplication_135 = multiplierReg_135 * io_man_b_135; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_7_T_17 = multiplication_135 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_135
    ; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_7_T_15 = {1'h0,dotProductRegs_2_7}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_7_T_16 = ~_two_complement_7_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_7_T_18 = _two_complement_7_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_136; // @[block_division.scala 204:34]
  reg  signReg_136; // @[block_division.scala 205:28]
  wire [9:0] multiplication_136 = multiplierReg_136 * io_man_b_136; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_8_T_17 = multiplication_136 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_136
    ; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_8_T_15 = {1'h0,dotProductRegs_2_8}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_8_T_16 = ~_two_complement_8_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_8_T_18 = _two_complement_8_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_137; // @[block_division.scala 204:34]
  reg  signReg_137; // @[block_division.scala 205:28]
  wire [9:0] multiplication_137 = multiplierReg_137 * io_man_b_137; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_9_T_17 = multiplication_137 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_137
    ; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_9_T_15 = {1'h0,dotProductRegs_2_9}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_9_T_16 = ~_two_complement_9_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_9_T_18 = _two_complement_9_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_138; // @[block_division.scala 204:34]
  reg  signReg_138; // @[block_division.scala 205:28]
  wire [9:0] multiplication_138 = multiplierReg_138 * io_man_b_138; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_10_T_17 = multiplication_138 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_138; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_10_T_15 = {1'h0,dotProductRegs_2_10}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_10_T_16 = ~_two_complement_10_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_10_T_18 = _two_complement_10_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_139; // @[block_division.scala 204:34]
  reg  signReg_139; // @[block_division.scala 205:28]
  wire [9:0] multiplication_139 = multiplierReg_139 * io_man_b_139; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_11_T_17 = multiplication_139 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_139; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_11_T_15 = {1'h0,dotProductRegs_2_11}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_11_T_16 = ~_two_complement_11_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_11_T_18 = _two_complement_11_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_140; // @[block_division.scala 204:34]
  reg  signReg_140; // @[block_division.scala 205:28]
  wire [9:0] multiplication_140 = multiplierReg_140 * io_man_b_140; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_12_T_17 = multiplication_140 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_140; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_12_T_15 = {1'h0,dotProductRegs_2_12}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_12_T_16 = ~_two_complement_12_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_12_T_18 = _two_complement_12_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_141; // @[block_division.scala 204:34]
  reg  signReg_141; // @[block_division.scala 205:28]
  wire [9:0] multiplication_141 = multiplierReg_141 * io_man_b_141; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_13_T_17 = multiplication_141 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_141; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_13_T_15 = {1'h0,dotProductRegs_2_13}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_13_T_16 = ~_two_complement_13_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_13_T_18 = _two_complement_13_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_142; // @[block_division.scala 204:34]
  reg  signReg_142; // @[block_division.scala 205:28]
  wire [9:0] multiplication_142 = multiplierReg_142 * io_man_b_142; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_14_T_17 = multiplication_142 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_142; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_14_T_15 = {1'h0,dotProductRegs_2_14}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_14_T_16 = ~_two_complement_14_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_14_T_18 = _two_complement_14_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_143; // @[block_division.scala 204:34]
  reg  signReg_143; // @[block_division.scala 205:28]
  wire [9:0] multiplication_143 = multiplierReg_143 * io_man_b_143; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_15_T_17 = multiplication_143 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_143; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_15_T_15 = {1'h0,dotProductRegs_2_15}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_15_T_16 = ~_two_complement_15_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_15_T_18 = _two_complement_15_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_144; // @[block_division.scala 204:34]
  reg  signReg_144; // @[block_division.scala 205:28]
  wire [9:0] multiplication_144 = multiplierReg_144 * io_man_b_144; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_16_T_17 = multiplication_144 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_144; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_16_T_15 = {1'h0,dotProductRegs_2_16}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_16_T_16 = ~_two_complement_16_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_16_T_18 = _two_complement_16_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_145; // @[block_division.scala 204:34]
  reg  signReg_145; // @[block_division.scala 205:28]
  wire [9:0] multiplication_145 = multiplierReg_145 * io_man_b_145; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_17_T_17 = multiplication_145 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_145; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_17_T_15 = {1'h0,dotProductRegs_2_17}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_17_T_16 = ~_two_complement_17_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_17_T_18 = _two_complement_17_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_146; // @[block_division.scala 204:34]
  reg  signReg_146; // @[block_division.scala 205:28]
  wire [9:0] multiplication_146 = multiplierReg_146 * io_man_b_146; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_18_T_17 = multiplication_146 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_146; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_18_T_15 = {1'h0,dotProductRegs_2_18}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_18_T_16 = ~_two_complement_18_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_18_T_18 = _two_complement_18_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_147; // @[block_division.scala 204:34]
  reg  signReg_147; // @[block_division.scala 205:28]
  wire [9:0] multiplication_147 = multiplierReg_147 * io_man_b_147; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_19_T_17 = multiplication_147 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_147; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_19_T_15 = {1'h0,dotProductRegs_2_19}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_19_T_16 = ~_two_complement_19_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_19_T_18 = _two_complement_19_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_148; // @[block_division.scala 204:34]
  reg  signReg_148; // @[block_division.scala 205:28]
  wire [9:0] multiplication_148 = multiplierReg_148 * io_man_b_148; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_20_T_17 = multiplication_148 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_148; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_20_T_15 = {1'h0,dotProductRegs_2_20}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_20_T_16 = ~_two_complement_20_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_20_T_18 = _two_complement_20_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_149; // @[block_division.scala 204:34]
  reg  signReg_149; // @[block_division.scala 205:28]
  wire [9:0] multiplication_149 = multiplierReg_149 * io_man_b_149; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_21_T_17 = multiplication_149 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_149; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_21_T_15 = {1'h0,dotProductRegs_2_21}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_21_T_16 = ~_two_complement_21_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_21_T_18 = _two_complement_21_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_150; // @[block_division.scala 204:34]
  reg  signReg_150; // @[block_division.scala 205:28]
  wire [9:0] multiplication_150 = multiplierReg_150 * io_man_b_150; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_22_T_17 = multiplication_150 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_150; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_22_T_15 = {1'h0,dotProductRegs_2_22}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_22_T_16 = ~_two_complement_22_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_22_T_18 = _two_complement_22_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_151; // @[block_division.scala 204:34]
  reg  signReg_151; // @[block_division.scala 205:28]
  wire [9:0] multiplication_151 = multiplierReg_151 * io_man_b_151; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_23_T_17 = multiplication_151 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_151; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_23_T_15 = {1'h0,dotProductRegs_2_23}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_23_T_16 = ~_two_complement_23_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_23_T_18 = _two_complement_23_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_152; // @[block_division.scala 204:34]
  reg  signReg_152; // @[block_division.scala 205:28]
  wire [9:0] multiplication_152 = multiplierReg_152 * io_man_b_152; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_24_T_17 = multiplication_152 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_152; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_24_T_15 = {1'h0,dotProductRegs_2_24}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_24_T_16 = ~_two_complement_24_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_24_T_18 = _two_complement_24_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_153; // @[block_division.scala 204:34]
  reg  signReg_153; // @[block_division.scala 205:28]
  wire [9:0] multiplication_153 = multiplierReg_153 * io_man_b_153; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_25_T_17 = multiplication_153 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_153; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_25_T_15 = {1'h0,dotProductRegs_2_25}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_25_T_16 = ~_two_complement_25_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_25_T_18 = _two_complement_25_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_154; // @[block_division.scala 204:34]
  reg  signReg_154; // @[block_division.scala 205:28]
  wire [9:0] multiplication_154 = multiplierReg_154 * io_man_b_154; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_26_T_17 = multiplication_154 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_154; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_26_T_15 = {1'h0,dotProductRegs_2_26}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_26_T_16 = ~_two_complement_26_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_26_T_18 = _two_complement_26_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_155; // @[block_division.scala 204:34]
  reg  signReg_155; // @[block_division.scala 205:28]
  wire [9:0] multiplication_155 = multiplierReg_155 * io_man_b_155; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_27_T_17 = multiplication_155 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_155; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_27_T_15 = {1'h0,dotProductRegs_2_27}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_27_T_16 = ~_two_complement_27_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_27_T_18 = _two_complement_27_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_156; // @[block_division.scala 204:34]
  reg  signReg_156; // @[block_division.scala 205:28]
  wire [9:0] multiplication_156 = multiplierReg_156 * io_man_b_156; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_28_T_17 = multiplication_156 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_156; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_28_T_15 = {1'h0,dotProductRegs_2_28}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_28_T_16 = ~_two_complement_28_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_28_T_18 = _two_complement_28_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_157; // @[block_division.scala 204:34]
  reg  signReg_157; // @[block_division.scala 205:28]
  wire [9:0] multiplication_157 = multiplierReg_157 * io_man_b_157; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_29_T_17 = multiplication_157 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_157; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_29_T_15 = {1'h0,dotProductRegs_2_29}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_29_T_16 = ~_two_complement_29_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_29_T_18 = _two_complement_29_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_158; // @[block_division.scala 204:34]
  reg  signReg_158; // @[block_division.scala 205:28]
  wire [9:0] multiplication_158 = multiplierReg_158 * io_man_b_158; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_30_T_17 = multiplication_158 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_158; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_30_T_15 = {1'h0,dotProductRegs_2_30}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_30_T_16 = ~_two_complement_30_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_30_T_18 = _two_complement_30_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_159; // @[block_division.scala 204:34]
  reg  signReg_159; // @[block_division.scala 205:28]
  wire [9:0] multiplication_159 = multiplierReg_159 * io_man_b_159; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_31_T_17 = multiplication_159 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_159; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_31_T_15 = {1'h0,dotProductRegs_2_31}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_31_T_16 = ~_two_complement_31_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_31_T_18 = _two_complement_31_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_160; // @[block_division.scala 204:34]
  reg  signReg_160; // @[block_division.scala 205:28]
  wire [9:0] multiplication_160 = multiplierReg_160 * io_man_b_160; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_32_T_17 = multiplication_160 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_160; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_32_T_15 = {1'h0,dotProductRegs_2_32}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_32_T_16 = ~_two_complement_32_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_32_T_18 = _two_complement_32_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_161; // @[block_division.scala 204:34]
  reg  signReg_161; // @[block_division.scala 205:28]
  wire [9:0] multiplication_161 = multiplierReg_161 * io_man_b_161; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_33_T_17 = multiplication_161 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_161; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_33_T_15 = {1'h0,dotProductRegs_2_33}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_33_T_16 = ~_two_complement_33_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_33_T_18 = _two_complement_33_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_162; // @[block_division.scala 204:34]
  reg  signReg_162; // @[block_division.scala 205:28]
  wire [9:0] multiplication_162 = multiplierReg_162 * io_man_b_162; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_34_T_17 = multiplication_162 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_162; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_34_T_15 = {1'h0,dotProductRegs_2_34}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_34_T_16 = ~_two_complement_34_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_34_T_18 = _two_complement_34_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_163; // @[block_division.scala 204:34]
  reg  signReg_163; // @[block_division.scala 205:28]
  wire [9:0] multiplication_163 = multiplierReg_163 * io_man_b_163; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_35_T_17 = multiplication_163 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_163; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_35_T_15 = {1'h0,dotProductRegs_2_35}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_35_T_16 = ~_two_complement_35_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_35_T_18 = _two_complement_35_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_164; // @[block_division.scala 204:34]
  reg  signReg_164; // @[block_division.scala 205:28]
  wire [9:0] multiplication_164 = multiplierReg_164 * io_man_b_164; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_36_T_17 = multiplication_164 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_164; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_36_T_15 = {1'h0,dotProductRegs_2_36}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_36_T_16 = ~_two_complement_36_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_36_T_18 = _two_complement_36_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_165; // @[block_division.scala 204:34]
  reg  signReg_165; // @[block_division.scala 205:28]
  wire [9:0] multiplication_165 = multiplierReg_165 * io_man_b_165; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_37_T_17 = multiplication_165 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_165; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_37_T_15 = {1'h0,dotProductRegs_2_37}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_37_T_16 = ~_two_complement_37_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_37_T_18 = _two_complement_37_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_166; // @[block_division.scala 204:34]
  reg  signReg_166; // @[block_division.scala 205:28]
  wire [9:0] multiplication_166 = multiplierReg_166 * io_man_b_166; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_38_T_17 = multiplication_166 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_166; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_38_T_15 = {1'h0,dotProductRegs_2_38}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_38_T_16 = ~_two_complement_38_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_38_T_18 = _two_complement_38_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_167; // @[block_division.scala 204:34]
  reg  signReg_167; // @[block_division.scala 205:28]
  wire [9:0] multiplication_167 = multiplierReg_167 * io_man_b_167; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_39_T_17 = multiplication_167 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_167; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_39_T_15 = {1'h0,dotProductRegs_2_39}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_39_T_16 = ~_two_complement_39_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_39_T_18 = _two_complement_39_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_168; // @[block_division.scala 204:34]
  reg  signReg_168; // @[block_division.scala 205:28]
  wire [9:0] multiplication_168 = multiplierReg_168 * io_man_b_168; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_40_T_17 = multiplication_168 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_168; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_40_T_15 = {1'h0,dotProductRegs_2_40}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_40_T_16 = ~_two_complement_40_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_40_T_18 = _two_complement_40_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_169; // @[block_division.scala 204:34]
  reg  signReg_169; // @[block_division.scala 205:28]
  wire [9:0] multiplication_169 = multiplierReg_169 * io_man_b_169; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_41_T_17 = multiplication_169 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_169; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_41_T_15 = {1'h0,dotProductRegs_2_41}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_41_T_16 = ~_two_complement_41_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_41_T_18 = _two_complement_41_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_170; // @[block_division.scala 204:34]
  reg  signReg_170; // @[block_division.scala 205:28]
  wire [9:0] multiplication_170 = multiplierReg_170 * io_man_b_170; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_42_T_17 = multiplication_170 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_170; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_42_T_15 = {1'h0,dotProductRegs_2_42}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_42_T_16 = ~_two_complement_42_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_42_T_18 = _two_complement_42_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_171; // @[block_division.scala 204:34]
  reg  signReg_171; // @[block_division.scala 205:28]
  wire [9:0] multiplication_171 = multiplierReg_171 * io_man_b_171; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_43_T_17 = multiplication_171 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_171; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_43_T_15 = {1'h0,dotProductRegs_2_43}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_43_T_16 = ~_two_complement_43_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_43_T_18 = _two_complement_43_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_172; // @[block_division.scala 204:34]
  reg  signReg_172; // @[block_division.scala 205:28]
  wire [9:0] multiplication_172 = multiplierReg_172 * io_man_b_172; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_44_T_17 = multiplication_172 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_172; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_44_T_15 = {1'h0,dotProductRegs_2_44}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_44_T_16 = ~_two_complement_44_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_44_T_18 = _two_complement_44_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_173; // @[block_division.scala 204:34]
  reg  signReg_173; // @[block_division.scala 205:28]
  wire [9:0] multiplication_173 = multiplierReg_173 * io_man_b_173; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_45_T_17 = multiplication_173 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_173; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_45_T_15 = {1'h0,dotProductRegs_2_45}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_45_T_16 = ~_two_complement_45_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_45_T_18 = _two_complement_45_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_174; // @[block_division.scala 204:34]
  reg  signReg_174; // @[block_division.scala 205:28]
  wire [9:0] multiplication_174 = multiplierReg_174 * io_man_b_174; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_46_T_17 = multiplication_174 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_174; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_46_T_15 = {1'h0,dotProductRegs_2_46}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_46_T_16 = ~_two_complement_46_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_46_T_18 = _two_complement_46_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_175; // @[block_division.scala 204:34]
  reg  signReg_175; // @[block_division.scala 205:28]
  wire [9:0] multiplication_175 = multiplierReg_175 * io_man_b_175; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_47_T_17 = multiplication_175 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_175; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_47_T_15 = {1'h0,dotProductRegs_2_47}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_47_T_16 = ~_two_complement_47_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_47_T_18 = _two_complement_47_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_176; // @[block_division.scala 204:34]
  reg  signReg_176; // @[block_division.scala 205:28]
  wire [9:0] multiplication_176 = multiplierReg_176 * io_man_b_176; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_48_T_17 = multiplication_176 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_176; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_48_T_15 = {1'h0,dotProductRegs_2_48}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_48_T_16 = ~_two_complement_48_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_48_T_18 = _two_complement_48_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_177; // @[block_division.scala 204:34]
  reg  signReg_177; // @[block_division.scala 205:28]
  wire [9:0] multiplication_177 = multiplierReg_177 * io_man_b_177; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_49_T_17 = multiplication_177 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_177; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_49_T_15 = {1'h0,dotProductRegs_2_49}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_49_T_16 = ~_two_complement_49_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_49_T_18 = _two_complement_49_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_178; // @[block_division.scala 204:34]
  reg  signReg_178; // @[block_division.scala 205:28]
  wire [9:0] multiplication_178 = multiplierReg_178 * io_man_b_178; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_50_T_17 = multiplication_178 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_178; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_50_T_15 = {1'h0,dotProductRegs_2_50}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_50_T_16 = ~_two_complement_50_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_50_T_18 = _two_complement_50_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_179; // @[block_division.scala 204:34]
  reg  signReg_179; // @[block_division.scala 205:28]
  wire [9:0] multiplication_179 = multiplierReg_179 * io_man_b_179; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_51_T_17 = multiplication_179 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_179; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_51_T_15 = {1'h0,dotProductRegs_2_51}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_51_T_16 = ~_two_complement_51_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_51_T_18 = _two_complement_51_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_180; // @[block_division.scala 204:34]
  reg  signReg_180; // @[block_division.scala 205:28]
  wire [9:0] multiplication_180 = multiplierReg_180 * io_man_b_180; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_52_T_17 = multiplication_180 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_180; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_52_T_15 = {1'h0,dotProductRegs_2_52}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_52_T_16 = ~_two_complement_52_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_52_T_18 = _two_complement_52_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_181; // @[block_division.scala 204:34]
  reg  signReg_181; // @[block_division.scala 205:28]
  wire [9:0] multiplication_181 = multiplierReg_181 * io_man_b_181; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_53_T_17 = multiplication_181 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_181; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_53_T_15 = {1'h0,dotProductRegs_2_53}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_53_T_16 = ~_two_complement_53_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_53_T_18 = _two_complement_53_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_182; // @[block_division.scala 204:34]
  reg  signReg_182; // @[block_division.scala 205:28]
  wire [9:0] multiplication_182 = multiplierReg_182 * io_man_b_182; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_54_T_17 = multiplication_182 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_182; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_54_T_15 = {1'h0,dotProductRegs_2_54}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_54_T_16 = ~_two_complement_54_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_54_T_18 = _two_complement_54_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_183; // @[block_division.scala 204:34]
  reg  signReg_183; // @[block_division.scala 205:28]
  wire [9:0] multiplication_183 = multiplierReg_183 * io_man_b_183; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_55_T_17 = multiplication_183 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_183; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_55_T_15 = {1'h0,dotProductRegs_2_55}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_55_T_16 = ~_two_complement_55_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_55_T_18 = _two_complement_55_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_184; // @[block_division.scala 204:34]
  reg  signReg_184; // @[block_division.scala 205:28]
  wire [9:0] multiplication_184 = multiplierReg_184 * io_man_b_184; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_56_T_17 = multiplication_184 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_184; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_56_T_15 = {1'h0,dotProductRegs_2_56}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_56_T_16 = ~_two_complement_56_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_56_T_18 = _two_complement_56_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_185; // @[block_division.scala 204:34]
  reg  signReg_185; // @[block_division.scala 205:28]
  wire [9:0] multiplication_185 = multiplierReg_185 * io_man_b_185; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_57_T_17 = multiplication_185 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_185; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_57_T_15 = {1'h0,dotProductRegs_2_57}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_57_T_16 = ~_two_complement_57_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_57_T_18 = _two_complement_57_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_186; // @[block_division.scala 204:34]
  reg  signReg_186; // @[block_division.scala 205:28]
  wire [9:0] multiplication_186 = multiplierReg_186 * io_man_b_186; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_58_T_17 = multiplication_186 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_186; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_58_T_15 = {1'h0,dotProductRegs_2_58}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_58_T_16 = ~_two_complement_58_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_58_T_18 = _two_complement_58_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_187; // @[block_division.scala 204:34]
  reg  signReg_187; // @[block_division.scala 205:28]
  wire [9:0] multiplication_187 = multiplierReg_187 * io_man_b_187; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_59_T_17 = multiplication_187 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_187; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_59_T_15 = {1'h0,dotProductRegs_2_59}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_59_T_16 = ~_two_complement_59_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_59_T_18 = _two_complement_59_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_188; // @[block_division.scala 204:34]
  reg  signReg_188; // @[block_division.scala 205:28]
  wire [9:0] multiplication_188 = multiplierReg_188 * io_man_b_188; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_60_T_17 = multiplication_188 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_188; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_60_T_15 = {1'h0,dotProductRegs_2_60}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_60_T_16 = ~_two_complement_60_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_60_T_18 = _two_complement_60_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_189; // @[block_division.scala 204:34]
  reg  signReg_189; // @[block_division.scala 205:28]
  wire [9:0] multiplication_189 = multiplierReg_189 * io_man_b_189; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_61_T_17 = multiplication_189 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_189; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_61_T_15 = {1'h0,dotProductRegs_2_61}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_61_T_16 = ~_two_complement_61_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_61_T_18 = _two_complement_61_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_190; // @[block_division.scala 204:34]
  reg  signReg_190; // @[block_division.scala 205:28]
  wire [9:0] multiplication_190 = multiplierReg_190 * io_man_b_190; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_62_T_17 = multiplication_190 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_190; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_62_T_15 = {1'h0,dotProductRegs_2_62}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_62_T_16 = ~_two_complement_62_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_62_T_18 = _two_complement_62_T_16 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_191; // @[block_division.scala 204:34]
  reg  signReg_191; // @[block_division.scala 205:28]
  wire [9:0] multiplication_191 = multiplierReg_191 * io_man_b_191; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_63_T_17 = multiplication_191 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_191; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_63_T_15 = {1'h0,dotProductRegs_2_63}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_63_T_16 = ~_two_complement_63_T_15; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_63_T_18 = _two_complement_63_T_16 + 6'h1; // @[block_division.scala 213:38]
  wire [6:0] _sum_T_124 = $signed(two_complement_buffer_2_0) + $signed(two_complement_buffer_2_1); // @[block_division.scala 218:46]
  wire [6:0] _GEN_320 = {{1{two_complement_buffer_2_2[5]}},two_complement_buffer_2_2}; // @[block_division.scala 218:46]
  wire [7:0] _sum_T_125 = $signed(_sum_T_124) + $signed(_GEN_320); // @[block_division.scala 218:46]
  wire [7:0] _GEN_321 = {{2{two_complement_buffer_2_3[5]}},two_complement_buffer_2_3}; // @[block_division.scala 218:46]
  wire [8:0] _sum_T_126 = $signed(_sum_T_125) + $signed(_GEN_321); // @[block_division.scala 218:46]
  wire [8:0] _GEN_322 = {{3{two_complement_buffer_2_4[5]}},two_complement_buffer_2_4}; // @[block_division.scala 218:46]
  wire [9:0] _sum_T_127 = $signed(_sum_T_126) + $signed(_GEN_322); // @[block_division.scala 218:46]
  wire [9:0] _GEN_323 = {{4{two_complement_buffer_2_5[5]}},two_complement_buffer_2_5}; // @[block_division.scala 218:46]
  wire [10:0] _sum_T_128 = $signed(_sum_T_127) + $signed(_GEN_323); // @[block_division.scala 218:46]
  wire [10:0] _GEN_324 = {{5{two_complement_buffer_2_6[5]}},two_complement_buffer_2_6}; // @[block_division.scala 218:46]
  wire [11:0] _sum_T_129 = $signed(_sum_T_128) + $signed(_GEN_324); // @[block_division.scala 218:46]
  wire [11:0] _GEN_325 = {{6{two_complement_buffer_2_7[5]}},two_complement_buffer_2_7}; // @[block_division.scala 218:46]
  wire [12:0] _sum_T_130 = $signed(_sum_T_129) + $signed(_GEN_325); // @[block_division.scala 218:46]
  wire [12:0] _GEN_326 = {{7{two_complement_buffer_2_8[5]}},two_complement_buffer_2_8}; // @[block_division.scala 218:46]
  wire [13:0] _sum_T_131 = $signed(_sum_T_130) + $signed(_GEN_326); // @[block_division.scala 218:46]
  wire [13:0] _GEN_327 = {{8{two_complement_buffer_2_9[5]}},two_complement_buffer_2_9}; // @[block_division.scala 218:46]
  wire [14:0] _sum_T_132 = $signed(_sum_T_131) + $signed(_GEN_327); // @[block_division.scala 218:46]
  wire [14:0] _GEN_328 = {{9{two_complement_buffer_2_10[5]}},two_complement_buffer_2_10}; // @[block_division.scala 218:46]
  wire [15:0] _sum_T_133 = $signed(_sum_T_132) + $signed(_GEN_328); // @[block_division.scala 218:46]
  wire [15:0] _GEN_329 = {{10{two_complement_buffer_2_11[5]}},two_complement_buffer_2_11}; // @[block_division.scala 218:46]
  wire [16:0] _sum_T_134 = $signed(_sum_T_133) + $signed(_GEN_329); // @[block_division.scala 218:46]
  wire [16:0] _GEN_330 = {{11{two_complement_buffer_2_12[5]}},two_complement_buffer_2_12}; // @[block_division.scala 218:46]
  wire [17:0] _sum_T_135 = $signed(_sum_T_134) + $signed(_GEN_330); // @[block_division.scala 218:46]
  wire [17:0] _GEN_331 = {{12{two_complement_buffer_2_13[5]}},two_complement_buffer_2_13}; // @[block_division.scala 218:46]
  wire [18:0] _sum_T_136 = $signed(_sum_T_135) + $signed(_GEN_331); // @[block_division.scala 218:46]
  wire [18:0] _GEN_332 = {{13{two_complement_buffer_2_14[5]}},two_complement_buffer_2_14}; // @[block_division.scala 218:46]
  wire [19:0] _sum_T_137 = $signed(_sum_T_136) + $signed(_GEN_332); // @[block_division.scala 218:46]
  wire [19:0] _GEN_333 = {{14{two_complement_buffer_2_15[5]}},two_complement_buffer_2_15}; // @[block_division.scala 218:46]
  wire [20:0] _sum_T_138 = $signed(_sum_T_137) + $signed(_GEN_333); // @[block_division.scala 218:46]
  wire [20:0] _GEN_334 = {{15{two_complement_buffer_2_16[5]}},two_complement_buffer_2_16}; // @[block_division.scala 218:46]
  wire [21:0] _sum_T_139 = $signed(_sum_T_138) + $signed(_GEN_334); // @[block_division.scala 218:46]
  wire [21:0] _GEN_335 = {{16{two_complement_buffer_2_17[5]}},two_complement_buffer_2_17}; // @[block_division.scala 218:46]
  wire [22:0] _sum_T_140 = $signed(_sum_T_139) + $signed(_GEN_335); // @[block_division.scala 218:46]
  wire [22:0] _GEN_336 = {{17{two_complement_buffer_2_18[5]}},two_complement_buffer_2_18}; // @[block_division.scala 218:46]
  wire [23:0] _sum_T_141 = $signed(_sum_T_140) + $signed(_GEN_336); // @[block_division.scala 218:46]
  wire [23:0] _GEN_337 = {{18{two_complement_buffer_2_19[5]}},two_complement_buffer_2_19}; // @[block_division.scala 218:46]
  wire [24:0] _sum_T_142 = $signed(_sum_T_141) + $signed(_GEN_337); // @[block_division.scala 218:46]
  wire [24:0] _GEN_338 = {{19{two_complement_buffer_2_20[5]}},two_complement_buffer_2_20}; // @[block_division.scala 218:46]
  wire [25:0] _sum_T_143 = $signed(_sum_T_142) + $signed(_GEN_338); // @[block_division.scala 218:46]
  wire [25:0] _GEN_339 = {{20{two_complement_buffer_2_21[5]}},two_complement_buffer_2_21}; // @[block_division.scala 218:46]
  wire [26:0] _sum_T_144 = $signed(_sum_T_143) + $signed(_GEN_339); // @[block_division.scala 218:46]
  wire [26:0] _GEN_340 = {{21{two_complement_buffer_2_22[5]}},two_complement_buffer_2_22}; // @[block_division.scala 218:46]
  wire [27:0] _sum_T_145 = $signed(_sum_T_144) + $signed(_GEN_340); // @[block_division.scala 218:46]
  wire [27:0] _GEN_341 = {{22{two_complement_buffer_2_23[5]}},two_complement_buffer_2_23}; // @[block_division.scala 218:46]
  wire [28:0] _sum_T_146 = $signed(_sum_T_145) + $signed(_GEN_341); // @[block_division.scala 218:46]
  wire [28:0] _GEN_342 = {{23{two_complement_buffer_2_24[5]}},two_complement_buffer_2_24}; // @[block_division.scala 218:46]
  wire [29:0] _sum_T_147 = $signed(_sum_T_146) + $signed(_GEN_342); // @[block_division.scala 218:46]
  wire [29:0] _GEN_343 = {{24{two_complement_buffer_2_25[5]}},two_complement_buffer_2_25}; // @[block_division.scala 218:46]
  wire [30:0] _sum_T_148 = $signed(_sum_T_147) + $signed(_GEN_343); // @[block_division.scala 218:46]
  wire [30:0] _GEN_344 = {{25{two_complement_buffer_2_26[5]}},two_complement_buffer_2_26}; // @[block_division.scala 218:46]
  wire [31:0] _sum_T_149 = $signed(_sum_T_148) + $signed(_GEN_344); // @[block_division.scala 218:46]
  wire [31:0] _GEN_345 = {{26{two_complement_buffer_2_27[5]}},two_complement_buffer_2_27}; // @[block_division.scala 218:46]
  wire [32:0] _sum_T_150 = $signed(_sum_T_149) + $signed(_GEN_345); // @[block_division.scala 218:46]
  wire [32:0] _GEN_346 = {{27{two_complement_buffer_2_28[5]}},two_complement_buffer_2_28}; // @[block_division.scala 218:46]
  wire [33:0] _sum_T_151 = $signed(_sum_T_150) + $signed(_GEN_346); // @[block_division.scala 218:46]
  wire [33:0] _GEN_347 = {{28{two_complement_buffer_2_29[5]}},two_complement_buffer_2_29}; // @[block_division.scala 218:46]
  wire [34:0] _sum_T_152 = $signed(_sum_T_151) + $signed(_GEN_347); // @[block_division.scala 218:46]
  wire [34:0] _GEN_348 = {{29{two_complement_buffer_2_30[5]}},two_complement_buffer_2_30}; // @[block_division.scala 218:46]
  wire [35:0] _sum_T_153 = $signed(_sum_T_152) + $signed(_GEN_348); // @[block_division.scala 218:46]
  wire [35:0] _GEN_349 = {{30{two_complement_buffer_2_31[5]}},two_complement_buffer_2_31}; // @[block_division.scala 218:46]
  wire [36:0] _sum_T_154 = $signed(_sum_T_153) + $signed(_GEN_349); // @[block_division.scala 218:46]
  wire [36:0] _GEN_350 = {{31{two_complement_buffer_2_32[5]}},two_complement_buffer_2_32}; // @[block_division.scala 218:46]
  wire [37:0] _sum_T_155 = $signed(_sum_T_154) + $signed(_GEN_350); // @[block_division.scala 218:46]
  wire [37:0] _GEN_351 = {{32{two_complement_buffer_2_33[5]}},two_complement_buffer_2_33}; // @[block_division.scala 218:46]
  wire [38:0] _sum_T_156 = $signed(_sum_T_155) + $signed(_GEN_351); // @[block_division.scala 218:46]
  wire [38:0] _GEN_352 = {{33{two_complement_buffer_2_34[5]}},two_complement_buffer_2_34}; // @[block_division.scala 218:46]
  wire [39:0] _sum_T_157 = $signed(_sum_T_156) + $signed(_GEN_352); // @[block_division.scala 218:46]
  wire [39:0] _GEN_353 = {{34{two_complement_buffer_2_35[5]}},two_complement_buffer_2_35}; // @[block_division.scala 218:46]
  wire [40:0] _sum_T_158 = $signed(_sum_T_157) + $signed(_GEN_353); // @[block_division.scala 218:46]
  wire [40:0] _GEN_354 = {{35{two_complement_buffer_2_36[5]}},two_complement_buffer_2_36}; // @[block_division.scala 218:46]
  wire [41:0] _sum_T_159 = $signed(_sum_T_158) + $signed(_GEN_354); // @[block_division.scala 218:46]
  wire [41:0] _GEN_355 = {{36{two_complement_buffer_2_37[5]}},two_complement_buffer_2_37}; // @[block_division.scala 218:46]
  wire [42:0] _sum_T_160 = $signed(_sum_T_159) + $signed(_GEN_355); // @[block_division.scala 218:46]
  wire [42:0] _GEN_356 = {{37{two_complement_buffer_2_38[5]}},two_complement_buffer_2_38}; // @[block_division.scala 218:46]
  wire [43:0] _sum_T_161 = $signed(_sum_T_160) + $signed(_GEN_356); // @[block_division.scala 218:46]
  wire [43:0] _GEN_357 = {{38{two_complement_buffer_2_39[5]}},two_complement_buffer_2_39}; // @[block_division.scala 218:46]
  wire [44:0] _sum_T_162 = $signed(_sum_T_161) + $signed(_GEN_357); // @[block_division.scala 218:46]
  wire [44:0] _GEN_358 = {{39{two_complement_buffer_2_40[5]}},two_complement_buffer_2_40}; // @[block_division.scala 218:46]
  wire [45:0] _sum_T_163 = $signed(_sum_T_162) + $signed(_GEN_358); // @[block_division.scala 218:46]
  wire [45:0] _GEN_359 = {{40{two_complement_buffer_2_41[5]}},two_complement_buffer_2_41}; // @[block_division.scala 218:46]
  wire [46:0] _sum_T_164 = $signed(_sum_T_163) + $signed(_GEN_359); // @[block_division.scala 218:46]
  wire [46:0] _GEN_360 = {{41{two_complement_buffer_2_42[5]}},two_complement_buffer_2_42}; // @[block_division.scala 218:46]
  wire [47:0] _sum_T_165 = $signed(_sum_T_164) + $signed(_GEN_360); // @[block_division.scala 218:46]
  wire [47:0] _GEN_361 = {{42{two_complement_buffer_2_43[5]}},two_complement_buffer_2_43}; // @[block_division.scala 218:46]
  wire [48:0] _sum_T_166 = $signed(_sum_T_165) + $signed(_GEN_361); // @[block_division.scala 218:46]
  wire [48:0] _GEN_362 = {{43{two_complement_buffer_2_44[5]}},two_complement_buffer_2_44}; // @[block_division.scala 218:46]
  wire [49:0] _sum_T_167 = $signed(_sum_T_166) + $signed(_GEN_362); // @[block_division.scala 218:46]
  wire [49:0] _GEN_363 = {{44{two_complement_buffer_2_45[5]}},two_complement_buffer_2_45}; // @[block_division.scala 218:46]
  wire [50:0] _sum_T_168 = $signed(_sum_T_167) + $signed(_GEN_363); // @[block_division.scala 218:46]
  wire [50:0] _GEN_364 = {{45{two_complement_buffer_2_46[5]}},two_complement_buffer_2_46}; // @[block_division.scala 218:46]
  wire [51:0] _sum_T_169 = $signed(_sum_T_168) + $signed(_GEN_364); // @[block_division.scala 218:46]
  wire [51:0] _GEN_365 = {{46{two_complement_buffer_2_47[5]}},two_complement_buffer_2_47}; // @[block_division.scala 218:46]
  wire [52:0] _sum_T_170 = $signed(_sum_T_169) + $signed(_GEN_365); // @[block_division.scala 218:46]
  wire [52:0] _GEN_366 = {{47{two_complement_buffer_2_48[5]}},two_complement_buffer_2_48}; // @[block_division.scala 218:46]
  wire [53:0] _sum_T_171 = $signed(_sum_T_170) + $signed(_GEN_366); // @[block_division.scala 218:46]
  wire [53:0] _GEN_367 = {{48{two_complement_buffer_2_49[5]}},two_complement_buffer_2_49}; // @[block_division.scala 218:46]
  wire [54:0] _sum_T_172 = $signed(_sum_T_171) + $signed(_GEN_367); // @[block_division.scala 218:46]
  wire [54:0] _GEN_368 = {{49{two_complement_buffer_2_50[5]}},two_complement_buffer_2_50}; // @[block_division.scala 218:46]
  wire [55:0] _sum_T_173 = $signed(_sum_T_172) + $signed(_GEN_368); // @[block_division.scala 218:46]
  wire [55:0] _GEN_369 = {{50{two_complement_buffer_2_51[5]}},two_complement_buffer_2_51}; // @[block_division.scala 218:46]
  wire [56:0] _sum_T_174 = $signed(_sum_T_173) + $signed(_GEN_369); // @[block_division.scala 218:46]
  wire [56:0] _GEN_370 = {{51{two_complement_buffer_2_52[5]}},two_complement_buffer_2_52}; // @[block_division.scala 218:46]
  wire [57:0] _sum_T_175 = $signed(_sum_T_174) + $signed(_GEN_370); // @[block_division.scala 218:46]
  wire [57:0] _GEN_371 = {{52{two_complement_buffer_2_53[5]}},two_complement_buffer_2_53}; // @[block_division.scala 218:46]
  wire [58:0] _sum_T_176 = $signed(_sum_T_175) + $signed(_GEN_371); // @[block_division.scala 218:46]
  wire [58:0] _GEN_372 = {{53{two_complement_buffer_2_54[5]}},two_complement_buffer_2_54}; // @[block_division.scala 218:46]
  wire [59:0] _sum_T_177 = $signed(_sum_T_176) + $signed(_GEN_372); // @[block_division.scala 218:46]
  wire [59:0] _GEN_373 = {{54{two_complement_buffer_2_55[5]}},two_complement_buffer_2_55}; // @[block_division.scala 218:46]
  wire [60:0] _sum_T_178 = $signed(_sum_T_177) + $signed(_GEN_373); // @[block_division.scala 218:46]
  wire [60:0] _GEN_374 = {{55{two_complement_buffer_2_56[5]}},two_complement_buffer_2_56}; // @[block_division.scala 218:46]
  wire [61:0] _sum_T_179 = $signed(_sum_T_178) + $signed(_GEN_374); // @[block_division.scala 218:46]
  wire [61:0] _GEN_375 = {{56{two_complement_buffer_2_57[5]}},two_complement_buffer_2_57}; // @[block_division.scala 218:46]
  wire [62:0] _sum_T_180 = $signed(_sum_T_179) + $signed(_GEN_375); // @[block_division.scala 218:46]
  wire [62:0] _GEN_376 = {{57{two_complement_buffer_2_58[5]}},two_complement_buffer_2_58}; // @[block_division.scala 218:46]
  wire [63:0] _sum_T_181 = $signed(_sum_T_180) + $signed(_GEN_376); // @[block_division.scala 218:46]
  wire [63:0] _GEN_377 = {{58{two_complement_buffer_2_59[5]}},two_complement_buffer_2_59}; // @[block_division.scala 218:46]
  wire [64:0] _sum_T_182 = $signed(_sum_T_181) + $signed(_GEN_377); // @[block_division.scala 218:46]
  wire [64:0] _GEN_378 = {{59{two_complement_buffer_2_60[5]}},two_complement_buffer_2_60}; // @[block_division.scala 218:46]
  wire [65:0] _sum_T_183 = $signed(_sum_T_182) + $signed(_GEN_378); // @[block_division.scala 218:46]
  wire [65:0] _GEN_379 = {{60{two_complement_buffer_2_61[5]}},two_complement_buffer_2_61}; // @[block_division.scala 218:46]
  wire [66:0] _sum_T_184 = $signed(_sum_T_183) + $signed(_GEN_379); // @[block_division.scala 218:46]
  wire [66:0] _GEN_380 = {{61{two_complement_buffer_2_62[5]}},two_complement_buffer_2_62}; // @[block_division.scala 218:46]
  wire [67:0] _sum_T_185 = $signed(_sum_T_184) + $signed(_GEN_380); // @[block_division.scala 218:46]
  wire [67:0] _GEN_381 = {{62{two_complement_buffer_2_63[5]}},two_complement_buffer_2_63}; // @[block_division.scala 218:46]
  wire [68:0] sum_2 = $signed(_sum_T_185) + $signed(_GEN_381); // @[block_division.scala 218:46]
  wire [67:0] _acc_2_T_3 = ~sum_2[67:0]; // @[block_division.scala 219:57]
  wire [67:0] _acc_2_T_5 = _acc_2_T_3 + 68'h1; // @[block_division.scala 219:86]
  wire [68:0] _acc_2_T_14 = $signed(_sum_T_185) + $signed(_GEN_381); // @[block_division.scala 219:145]
  wire [68:0] _acc_2_T_15 = _acc_2_T_5 > _GEN_126 ? {{63'd0}, _acc_0_T_13} : _acc_2_T_14; // @[block_division.scala 219:55]
  wire [68:0] _acc_2_T_23 = sum_2[67:0] > _GEN_126 ? {{63'd0}, _dotProductRegs_0_T_1} : _acc_2_T_14; // @[block_division.scala 220:6]
  wire [68:0] _acc_2_T_24 = sum_2[68] ? _acc_2_T_15 : _acc_2_T_23; // @[block_division.scala 219:18]
  wire [8:0] _exp_output_3_T = io_exp_a_3 + io_exp_b_3; // @[block_division.scala 198:34]
  reg [4:0] dotProductRegs_3_0; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_1; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_2; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_3; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_4; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_5; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_6; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_7; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_8; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_9; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_10; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_11; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_12; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_13; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_14; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_15; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_16; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_17; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_18; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_19; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_20; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_21; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_22; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_23; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_24; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_25; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_26; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_27; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_28; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_29; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_30; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_31; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_32; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_33; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_34; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_35; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_36; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_37; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_38; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_39; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_40; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_41; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_42; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_43; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_44; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_45; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_46; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_47; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_48; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_49; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_50; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_51; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_52; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_53; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_54; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_55; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_56; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_57; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_58; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_59; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_60; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_61; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_62; // @[block_division.scala 199:29]
  reg [4:0] dotProductRegs_3_63; // @[block_division.scala 199:29]
  reg  signs_3_0; // @[block_division.scala 200:20]
  reg  signs_3_1; // @[block_division.scala 200:20]
  reg  signs_3_2; // @[block_division.scala 200:20]
  reg  signs_3_3; // @[block_division.scala 200:20]
  reg  signs_3_4; // @[block_division.scala 200:20]
  reg  signs_3_5; // @[block_division.scala 200:20]
  reg  signs_3_6; // @[block_division.scala 200:20]
  reg  signs_3_7; // @[block_division.scala 200:20]
  reg  signs_3_8; // @[block_division.scala 200:20]
  reg  signs_3_9; // @[block_division.scala 200:20]
  reg  signs_3_10; // @[block_division.scala 200:20]
  reg  signs_3_11; // @[block_division.scala 200:20]
  reg  signs_3_12; // @[block_division.scala 200:20]
  reg  signs_3_13; // @[block_division.scala 200:20]
  reg  signs_3_14; // @[block_division.scala 200:20]
  reg  signs_3_15; // @[block_division.scala 200:20]
  reg  signs_3_16; // @[block_division.scala 200:20]
  reg  signs_3_17; // @[block_division.scala 200:20]
  reg  signs_3_18; // @[block_division.scala 200:20]
  reg  signs_3_19; // @[block_division.scala 200:20]
  reg  signs_3_20; // @[block_division.scala 200:20]
  reg  signs_3_21; // @[block_division.scala 200:20]
  reg  signs_3_22; // @[block_division.scala 200:20]
  reg  signs_3_23; // @[block_division.scala 200:20]
  reg  signs_3_24; // @[block_division.scala 200:20]
  reg  signs_3_25; // @[block_division.scala 200:20]
  reg  signs_3_26; // @[block_division.scala 200:20]
  reg  signs_3_27; // @[block_division.scala 200:20]
  reg  signs_3_28; // @[block_division.scala 200:20]
  reg  signs_3_29; // @[block_division.scala 200:20]
  reg  signs_3_30; // @[block_division.scala 200:20]
  reg  signs_3_31; // @[block_division.scala 200:20]
  reg  signs_3_32; // @[block_division.scala 200:20]
  reg  signs_3_33; // @[block_division.scala 200:20]
  reg  signs_3_34; // @[block_division.scala 200:20]
  reg  signs_3_35; // @[block_division.scala 200:20]
  reg  signs_3_36; // @[block_division.scala 200:20]
  reg  signs_3_37; // @[block_division.scala 200:20]
  reg  signs_3_38; // @[block_division.scala 200:20]
  reg  signs_3_39; // @[block_division.scala 200:20]
  reg  signs_3_40; // @[block_division.scala 200:20]
  reg  signs_3_41; // @[block_division.scala 200:20]
  reg  signs_3_42; // @[block_division.scala 200:20]
  reg  signs_3_43; // @[block_division.scala 200:20]
  reg  signs_3_44; // @[block_division.scala 200:20]
  reg  signs_3_45; // @[block_division.scala 200:20]
  reg  signs_3_46; // @[block_division.scala 200:20]
  reg  signs_3_47; // @[block_division.scala 200:20]
  reg  signs_3_48; // @[block_division.scala 200:20]
  reg  signs_3_49; // @[block_division.scala 200:20]
  reg  signs_3_50; // @[block_division.scala 200:20]
  reg  signs_3_51; // @[block_division.scala 200:20]
  reg  signs_3_52; // @[block_division.scala 200:20]
  reg  signs_3_53; // @[block_division.scala 200:20]
  reg  signs_3_54; // @[block_division.scala 200:20]
  reg  signs_3_55; // @[block_division.scala 200:20]
  reg  signs_3_56; // @[block_division.scala 200:20]
  reg  signs_3_57; // @[block_division.scala 200:20]
  reg  signs_3_58; // @[block_division.scala 200:20]
  reg  signs_3_59; // @[block_division.scala 200:20]
  reg  signs_3_60; // @[block_division.scala 200:20]
  reg  signs_3_61; // @[block_division.scala 200:20]
  reg  signs_3_62; // @[block_division.scala 200:20]
  reg  signs_3_63; // @[block_division.scala 200:20]
  reg [5:0] two_complement_3_0; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_1; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_2; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_3; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_4; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_5; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_6; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_7; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_8; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_9; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_10; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_11; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_12; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_13; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_14; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_15; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_16; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_17; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_18; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_19; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_20; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_21; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_22; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_23; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_24; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_25; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_26; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_27; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_28; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_29; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_30; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_31; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_32; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_33; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_34; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_35; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_36; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_37; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_38; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_39; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_40; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_41; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_42; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_43; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_44; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_45; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_46; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_47; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_48; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_49; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_50; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_51; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_52; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_53; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_54; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_55; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_56; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_57; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_58; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_59; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_60; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_61; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_62; // @[block_division.scala 201:29]
  reg [5:0] two_complement_3_63; // @[block_division.scala 201:29]
  reg [5:0] two_complement_buffer_3_0; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_1; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_2; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_3; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_4; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_5; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_6; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_7; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_8; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_9; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_10; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_11; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_12; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_13; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_14; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_15; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_16; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_17; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_18; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_19; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_20; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_21; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_22; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_23; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_24; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_25; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_26; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_27; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_28; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_29; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_30; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_31; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_32; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_33; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_34; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_35; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_36; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_37; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_38; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_39; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_40; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_41; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_42; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_43; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_44; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_45; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_46; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_47; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_48; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_49; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_50; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_51; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_52; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_53; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_54; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_55; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_56; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_57; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_58; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_59; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_60; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_61; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_62; // @[block_division.scala 202:36]
  reg [5:0] two_complement_buffer_3_63; // @[block_division.scala 202:36]
  reg [4:0] multiplierReg_192; // @[block_division.scala 204:34]
  reg  signReg_192; // @[block_division.scala 205:28]
  wire [9:0] multiplication_192 = multiplierReg_192 * io_man_b_192; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_0_T_23 = multiplication_192 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_192
    ; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_0_T_22 = {1'h0,dotProductRegs_3_0}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_0_T_23 = ~_two_complement_0_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_0_T_25 = _two_complement_0_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_193; // @[block_division.scala 204:34]
  reg  signReg_193; // @[block_division.scala 205:28]
  wire [9:0] multiplication_193 = multiplierReg_193 * io_man_b_193; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_1_T_23 = multiplication_193 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_193
    ; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_1_T_22 = {1'h0,dotProductRegs_3_1}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_1_T_23 = ~_two_complement_1_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_1_T_25 = _two_complement_1_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_194; // @[block_division.scala 204:34]
  reg  signReg_194; // @[block_division.scala 205:28]
  wire [9:0] multiplication_194 = multiplierReg_194 * io_man_b_194; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_2_T_23 = multiplication_194 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_194
    ; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_2_T_22 = {1'h0,dotProductRegs_3_2}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_2_T_23 = ~_two_complement_2_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_2_T_25 = _two_complement_2_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_195; // @[block_division.scala 204:34]
  reg  signReg_195; // @[block_division.scala 205:28]
  wire [9:0] multiplication_195 = multiplierReg_195 * io_man_b_195; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_3_T_23 = multiplication_195 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_195
    ; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_3_T_22 = {1'h0,dotProductRegs_3_3}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_3_T_23 = ~_two_complement_3_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_3_T_25 = _two_complement_3_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_196; // @[block_division.scala 204:34]
  reg  signReg_196; // @[block_division.scala 205:28]
  wire [9:0] multiplication_196 = multiplierReg_196 * io_man_b_196; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_4_T_23 = multiplication_196 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_196
    ; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_4_T_22 = {1'h0,dotProductRegs_3_4}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_4_T_23 = ~_two_complement_4_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_4_T_25 = _two_complement_4_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_197; // @[block_division.scala 204:34]
  reg  signReg_197; // @[block_division.scala 205:28]
  wire [9:0] multiplication_197 = multiplierReg_197 * io_man_b_197; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_5_T_23 = multiplication_197 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_197
    ; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_5_T_22 = {1'h0,dotProductRegs_3_5}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_5_T_23 = ~_two_complement_5_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_5_T_25 = _two_complement_5_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_198; // @[block_division.scala 204:34]
  reg  signReg_198; // @[block_division.scala 205:28]
  wire [9:0] multiplication_198 = multiplierReg_198 * io_man_b_198; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_6_T_23 = multiplication_198 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_198
    ; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_6_T_22 = {1'h0,dotProductRegs_3_6}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_6_T_23 = ~_two_complement_6_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_6_T_25 = _two_complement_6_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_199; // @[block_division.scala 204:34]
  reg  signReg_199; // @[block_division.scala 205:28]
  wire [9:0] multiplication_199 = multiplierReg_199 * io_man_b_199; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_7_T_23 = multiplication_199 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_199
    ; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_7_T_22 = {1'h0,dotProductRegs_3_7}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_7_T_23 = ~_two_complement_7_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_7_T_25 = _two_complement_7_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_200; // @[block_division.scala 204:34]
  reg  signReg_200; // @[block_division.scala 205:28]
  wire [9:0] multiplication_200 = multiplierReg_200 * io_man_b_200; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_8_T_23 = multiplication_200 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_200
    ; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_8_T_22 = {1'h0,dotProductRegs_3_8}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_8_T_23 = ~_two_complement_8_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_8_T_25 = _two_complement_8_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_201; // @[block_division.scala 204:34]
  reg  signReg_201; // @[block_division.scala 205:28]
  wire [9:0] multiplication_201 = multiplierReg_201 * io_man_b_201; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_9_T_23 = multiplication_201 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} : multiplication_201
    ; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_9_T_22 = {1'h0,dotProductRegs_3_9}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_9_T_23 = ~_two_complement_9_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_9_T_25 = _two_complement_9_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_202; // @[block_division.scala 204:34]
  reg  signReg_202; // @[block_division.scala 205:28]
  wire [9:0] multiplication_202 = multiplierReg_202 * io_man_b_202; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_10_T_23 = multiplication_202 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_202; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_10_T_22 = {1'h0,dotProductRegs_3_10}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_10_T_23 = ~_two_complement_10_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_10_T_25 = _two_complement_10_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_203; // @[block_division.scala 204:34]
  reg  signReg_203; // @[block_division.scala 205:28]
  wire [9:0] multiplication_203 = multiplierReg_203 * io_man_b_203; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_11_T_23 = multiplication_203 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_203; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_11_T_22 = {1'h0,dotProductRegs_3_11}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_11_T_23 = ~_two_complement_11_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_11_T_25 = _two_complement_11_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_204; // @[block_division.scala 204:34]
  reg  signReg_204; // @[block_division.scala 205:28]
  wire [9:0] multiplication_204 = multiplierReg_204 * io_man_b_204; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_12_T_23 = multiplication_204 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_204; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_12_T_22 = {1'h0,dotProductRegs_3_12}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_12_T_23 = ~_two_complement_12_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_12_T_25 = _two_complement_12_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_205; // @[block_division.scala 204:34]
  reg  signReg_205; // @[block_division.scala 205:28]
  wire [9:0] multiplication_205 = multiplierReg_205 * io_man_b_205; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_13_T_23 = multiplication_205 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_205; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_13_T_22 = {1'h0,dotProductRegs_3_13}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_13_T_23 = ~_two_complement_13_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_13_T_25 = _two_complement_13_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_206; // @[block_division.scala 204:34]
  reg  signReg_206; // @[block_division.scala 205:28]
  wire [9:0] multiplication_206 = multiplierReg_206 * io_man_b_206; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_14_T_23 = multiplication_206 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_206; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_14_T_22 = {1'h0,dotProductRegs_3_14}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_14_T_23 = ~_two_complement_14_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_14_T_25 = _two_complement_14_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_207; // @[block_division.scala 204:34]
  reg  signReg_207; // @[block_division.scala 205:28]
  wire [9:0] multiplication_207 = multiplierReg_207 * io_man_b_207; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_15_T_23 = multiplication_207 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_207; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_15_T_22 = {1'h0,dotProductRegs_3_15}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_15_T_23 = ~_two_complement_15_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_15_T_25 = _two_complement_15_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_208; // @[block_division.scala 204:34]
  reg  signReg_208; // @[block_division.scala 205:28]
  wire [9:0] multiplication_208 = multiplierReg_208 * io_man_b_208; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_16_T_23 = multiplication_208 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_208; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_16_T_22 = {1'h0,dotProductRegs_3_16}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_16_T_23 = ~_two_complement_16_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_16_T_25 = _two_complement_16_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_209; // @[block_division.scala 204:34]
  reg  signReg_209; // @[block_division.scala 205:28]
  wire [9:0] multiplication_209 = multiplierReg_209 * io_man_b_209; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_17_T_23 = multiplication_209 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_209; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_17_T_22 = {1'h0,dotProductRegs_3_17}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_17_T_23 = ~_two_complement_17_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_17_T_25 = _two_complement_17_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_210; // @[block_division.scala 204:34]
  reg  signReg_210; // @[block_division.scala 205:28]
  wire [9:0] multiplication_210 = multiplierReg_210 * io_man_b_210; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_18_T_23 = multiplication_210 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_210; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_18_T_22 = {1'h0,dotProductRegs_3_18}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_18_T_23 = ~_two_complement_18_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_18_T_25 = _two_complement_18_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_211; // @[block_division.scala 204:34]
  reg  signReg_211; // @[block_division.scala 205:28]
  wire [9:0] multiplication_211 = multiplierReg_211 * io_man_b_211; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_19_T_23 = multiplication_211 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_211; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_19_T_22 = {1'h0,dotProductRegs_3_19}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_19_T_23 = ~_two_complement_19_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_19_T_25 = _two_complement_19_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_212; // @[block_division.scala 204:34]
  reg  signReg_212; // @[block_division.scala 205:28]
  wire [9:0] multiplication_212 = multiplierReg_212 * io_man_b_212; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_20_T_23 = multiplication_212 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_212; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_20_T_22 = {1'h0,dotProductRegs_3_20}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_20_T_23 = ~_two_complement_20_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_20_T_25 = _two_complement_20_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_213; // @[block_division.scala 204:34]
  reg  signReg_213; // @[block_division.scala 205:28]
  wire [9:0] multiplication_213 = multiplierReg_213 * io_man_b_213; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_21_T_23 = multiplication_213 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_213; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_21_T_22 = {1'h0,dotProductRegs_3_21}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_21_T_23 = ~_two_complement_21_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_21_T_25 = _two_complement_21_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_214; // @[block_division.scala 204:34]
  reg  signReg_214; // @[block_division.scala 205:28]
  wire [9:0] multiplication_214 = multiplierReg_214 * io_man_b_214; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_22_T_23 = multiplication_214 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_214; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_22_T_22 = {1'h0,dotProductRegs_3_22}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_22_T_23 = ~_two_complement_22_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_22_T_25 = _two_complement_22_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_215; // @[block_division.scala 204:34]
  reg  signReg_215; // @[block_division.scala 205:28]
  wire [9:0] multiplication_215 = multiplierReg_215 * io_man_b_215; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_23_T_23 = multiplication_215 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_215; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_23_T_22 = {1'h0,dotProductRegs_3_23}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_23_T_23 = ~_two_complement_23_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_23_T_25 = _two_complement_23_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_216; // @[block_division.scala 204:34]
  reg  signReg_216; // @[block_division.scala 205:28]
  wire [9:0] multiplication_216 = multiplierReg_216 * io_man_b_216; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_24_T_23 = multiplication_216 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_216; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_24_T_22 = {1'h0,dotProductRegs_3_24}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_24_T_23 = ~_two_complement_24_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_24_T_25 = _two_complement_24_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_217; // @[block_division.scala 204:34]
  reg  signReg_217; // @[block_division.scala 205:28]
  wire [9:0] multiplication_217 = multiplierReg_217 * io_man_b_217; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_25_T_23 = multiplication_217 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_217; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_25_T_22 = {1'h0,dotProductRegs_3_25}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_25_T_23 = ~_two_complement_25_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_25_T_25 = _two_complement_25_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_218; // @[block_division.scala 204:34]
  reg  signReg_218; // @[block_division.scala 205:28]
  wire [9:0] multiplication_218 = multiplierReg_218 * io_man_b_218; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_26_T_23 = multiplication_218 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_218; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_26_T_22 = {1'h0,dotProductRegs_3_26}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_26_T_23 = ~_two_complement_26_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_26_T_25 = _two_complement_26_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_219; // @[block_division.scala 204:34]
  reg  signReg_219; // @[block_division.scala 205:28]
  wire [9:0] multiplication_219 = multiplierReg_219 * io_man_b_219; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_27_T_23 = multiplication_219 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_219; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_27_T_22 = {1'h0,dotProductRegs_3_27}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_27_T_23 = ~_two_complement_27_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_27_T_25 = _two_complement_27_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_220; // @[block_division.scala 204:34]
  reg  signReg_220; // @[block_division.scala 205:28]
  wire [9:0] multiplication_220 = multiplierReg_220 * io_man_b_220; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_28_T_23 = multiplication_220 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_220; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_28_T_22 = {1'h0,dotProductRegs_3_28}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_28_T_23 = ~_two_complement_28_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_28_T_25 = _two_complement_28_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_221; // @[block_division.scala 204:34]
  reg  signReg_221; // @[block_division.scala 205:28]
  wire [9:0] multiplication_221 = multiplierReg_221 * io_man_b_221; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_29_T_23 = multiplication_221 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_221; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_29_T_22 = {1'h0,dotProductRegs_3_29}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_29_T_23 = ~_two_complement_29_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_29_T_25 = _two_complement_29_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_222; // @[block_division.scala 204:34]
  reg  signReg_222; // @[block_division.scala 205:28]
  wire [9:0] multiplication_222 = multiplierReg_222 * io_man_b_222; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_30_T_23 = multiplication_222 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_222; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_30_T_22 = {1'h0,dotProductRegs_3_30}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_30_T_23 = ~_two_complement_30_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_30_T_25 = _two_complement_30_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_223; // @[block_division.scala 204:34]
  reg  signReg_223; // @[block_division.scala 205:28]
  wire [9:0] multiplication_223 = multiplierReg_223 * io_man_b_223; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_31_T_23 = multiplication_223 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_223; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_31_T_22 = {1'h0,dotProductRegs_3_31}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_31_T_23 = ~_two_complement_31_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_31_T_25 = _two_complement_31_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_224; // @[block_division.scala 204:34]
  reg  signReg_224; // @[block_division.scala 205:28]
  wire [9:0] multiplication_224 = multiplierReg_224 * io_man_b_224; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_32_T_23 = multiplication_224 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_224; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_32_T_22 = {1'h0,dotProductRegs_3_32}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_32_T_23 = ~_two_complement_32_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_32_T_25 = _two_complement_32_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_225; // @[block_division.scala 204:34]
  reg  signReg_225; // @[block_division.scala 205:28]
  wire [9:0] multiplication_225 = multiplierReg_225 * io_man_b_225; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_33_T_23 = multiplication_225 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_225; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_33_T_22 = {1'h0,dotProductRegs_3_33}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_33_T_23 = ~_two_complement_33_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_33_T_25 = _two_complement_33_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_226; // @[block_division.scala 204:34]
  reg  signReg_226; // @[block_division.scala 205:28]
  wire [9:0] multiplication_226 = multiplierReg_226 * io_man_b_226; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_34_T_23 = multiplication_226 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_226; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_34_T_22 = {1'h0,dotProductRegs_3_34}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_34_T_23 = ~_two_complement_34_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_34_T_25 = _two_complement_34_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_227; // @[block_division.scala 204:34]
  reg  signReg_227; // @[block_division.scala 205:28]
  wire [9:0] multiplication_227 = multiplierReg_227 * io_man_b_227; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_35_T_23 = multiplication_227 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_227; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_35_T_22 = {1'h0,dotProductRegs_3_35}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_35_T_23 = ~_two_complement_35_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_35_T_25 = _two_complement_35_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_228; // @[block_division.scala 204:34]
  reg  signReg_228; // @[block_division.scala 205:28]
  wire [9:0] multiplication_228 = multiplierReg_228 * io_man_b_228; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_36_T_23 = multiplication_228 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_228; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_36_T_22 = {1'h0,dotProductRegs_3_36}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_36_T_23 = ~_two_complement_36_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_36_T_25 = _two_complement_36_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_229; // @[block_division.scala 204:34]
  reg  signReg_229; // @[block_division.scala 205:28]
  wire [9:0] multiplication_229 = multiplierReg_229 * io_man_b_229; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_37_T_23 = multiplication_229 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_229; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_37_T_22 = {1'h0,dotProductRegs_3_37}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_37_T_23 = ~_two_complement_37_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_37_T_25 = _two_complement_37_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_230; // @[block_division.scala 204:34]
  reg  signReg_230; // @[block_division.scala 205:28]
  wire [9:0] multiplication_230 = multiplierReg_230 * io_man_b_230; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_38_T_23 = multiplication_230 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_230; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_38_T_22 = {1'h0,dotProductRegs_3_38}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_38_T_23 = ~_two_complement_38_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_38_T_25 = _two_complement_38_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_231; // @[block_division.scala 204:34]
  reg  signReg_231; // @[block_division.scala 205:28]
  wire [9:0] multiplication_231 = multiplierReg_231 * io_man_b_231; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_39_T_23 = multiplication_231 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_231; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_39_T_22 = {1'h0,dotProductRegs_3_39}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_39_T_23 = ~_two_complement_39_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_39_T_25 = _two_complement_39_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_232; // @[block_division.scala 204:34]
  reg  signReg_232; // @[block_division.scala 205:28]
  wire [9:0] multiplication_232 = multiplierReg_232 * io_man_b_232; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_40_T_23 = multiplication_232 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_232; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_40_T_22 = {1'h0,dotProductRegs_3_40}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_40_T_23 = ~_two_complement_40_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_40_T_25 = _two_complement_40_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_233; // @[block_division.scala 204:34]
  reg  signReg_233; // @[block_division.scala 205:28]
  wire [9:0] multiplication_233 = multiplierReg_233 * io_man_b_233; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_41_T_23 = multiplication_233 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_233; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_41_T_22 = {1'h0,dotProductRegs_3_41}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_41_T_23 = ~_two_complement_41_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_41_T_25 = _two_complement_41_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_234; // @[block_division.scala 204:34]
  reg  signReg_234; // @[block_division.scala 205:28]
  wire [9:0] multiplication_234 = multiplierReg_234 * io_man_b_234; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_42_T_23 = multiplication_234 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_234; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_42_T_22 = {1'h0,dotProductRegs_3_42}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_42_T_23 = ~_two_complement_42_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_42_T_25 = _two_complement_42_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_235; // @[block_division.scala 204:34]
  reg  signReg_235; // @[block_division.scala 205:28]
  wire [9:0] multiplication_235 = multiplierReg_235 * io_man_b_235; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_43_T_23 = multiplication_235 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_235; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_43_T_22 = {1'h0,dotProductRegs_3_43}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_43_T_23 = ~_two_complement_43_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_43_T_25 = _two_complement_43_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_236; // @[block_division.scala 204:34]
  reg  signReg_236; // @[block_division.scala 205:28]
  wire [9:0] multiplication_236 = multiplierReg_236 * io_man_b_236; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_44_T_23 = multiplication_236 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_236; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_44_T_22 = {1'h0,dotProductRegs_3_44}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_44_T_23 = ~_two_complement_44_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_44_T_25 = _two_complement_44_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_237; // @[block_division.scala 204:34]
  reg  signReg_237; // @[block_division.scala 205:28]
  wire [9:0] multiplication_237 = multiplierReg_237 * io_man_b_237; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_45_T_23 = multiplication_237 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_237; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_45_T_22 = {1'h0,dotProductRegs_3_45}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_45_T_23 = ~_two_complement_45_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_45_T_25 = _two_complement_45_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_238; // @[block_division.scala 204:34]
  reg  signReg_238; // @[block_division.scala 205:28]
  wire [9:0] multiplication_238 = multiplierReg_238 * io_man_b_238; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_46_T_23 = multiplication_238 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_238; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_46_T_22 = {1'h0,dotProductRegs_3_46}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_46_T_23 = ~_two_complement_46_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_46_T_25 = _two_complement_46_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_239; // @[block_division.scala 204:34]
  reg  signReg_239; // @[block_division.scala 205:28]
  wire [9:0] multiplication_239 = multiplierReg_239 * io_man_b_239; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_47_T_23 = multiplication_239 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_239; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_47_T_22 = {1'h0,dotProductRegs_3_47}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_47_T_23 = ~_two_complement_47_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_47_T_25 = _two_complement_47_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_240; // @[block_division.scala 204:34]
  reg  signReg_240; // @[block_division.scala 205:28]
  wire [9:0] multiplication_240 = multiplierReg_240 * io_man_b_240; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_48_T_23 = multiplication_240 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_240; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_48_T_22 = {1'h0,dotProductRegs_3_48}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_48_T_23 = ~_two_complement_48_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_48_T_25 = _two_complement_48_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_241; // @[block_division.scala 204:34]
  reg  signReg_241; // @[block_division.scala 205:28]
  wire [9:0] multiplication_241 = multiplierReg_241 * io_man_b_241; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_49_T_23 = multiplication_241 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_241; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_49_T_22 = {1'h0,dotProductRegs_3_49}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_49_T_23 = ~_two_complement_49_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_49_T_25 = _two_complement_49_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_242; // @[block_division.scala 204:34]
  reg  signReg_242; // @[block_division.scala 205:28]
  wire [9:0] multiplication_242 = multiplierReg_242 * io_man_b_242; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_50_T_23 = multiplication_242 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_242; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_50_T_22 = {1'h0,dotProductRegs_3_50}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_50_T_23 = ~_two_complement_50_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_50_T_25 = _two_complement_50_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_243; // @[block_division.scala 204:34]
  reg  signReg_243; // @[block_division.scala 205:28]
  wire [9:0] multiplication_243 = multiplierReg_243 * io_man_b_243; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_51_T_23 = multiplication_243 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_243; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_51_T_22 = {1'h0,dotProductRegs_3_51}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_51_T_23 = ~_two_complement_51_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_51_T_25 = _two_complement_51_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_244; // @[block_division.scala 204:34]
  reg  signReg_244; // @[block_division.scala 205:28]
  wire [9:0] multiplication_244 = multiplierReg_244 * io_man_b_244; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_52_T_23 = multiplication_244 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_244; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_52_T_22 = {1'h0,dotProductRegs_3_52}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_52_T_23 = ~_two_complement_52_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_52_T_25 = _two_complement_52_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_245; // @[block_division.scala 204:34]
  reg  signReg_245; // @[block_division.scala 205:28]
  wire [9:0] multiplication_245 = multiplierReg_245 * io_man_b_245; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_53_T_23 = multiplication_245 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_245; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_53_T_22 = {1'h0,dotProductRegs_3_53}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_53_T_23 = ~_two_complement_53_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_53_T_25 = _two_complement_53_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_246; // @[block_division.scala 204:34]
  reg  signReg_246; // @[block_division.scala 205:28]
  wire [9:0] multiplication_246 = multiplierReg_246 * io_man_b_246; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_54_T_23 = multiplication_246 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_246; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_54_T_22 = {1'h0,dotProductRegs_3_54}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_54_T_23 = ~_two_complement_54_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_54_T_25 = _two_complement_54_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_247; // @[block_division.scala 204:34]
  reg  signReg_247; // @[block_division.scala 205:28]
  wire [9:0] multiplication_247 = multiplierReg_247 * io_man_b_247; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_55_T_23 = multiplication_247 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_247; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_55_T_22 = {1'h0,dotProductRegs_3_55}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_55_T_23 = ~_two_complement_55_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_55_T_25 = _two_complement_55_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_248; // @[block_division.scala 204:34]
  reg  signReg_248; // @[block_division.scala 205:28]
  wire [9:0] multiplication_248 = multiplierReg_248 * io_man_b_248; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_56_T_23 = multiplication_248 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_248; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_56_T_22 = {1'h0,dotProductRegs_3_56}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_56_T_23 = ~_two_complement_56_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_56_T_25 = _two_complement_56_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_249; // @[block_division.scala 204:34]
  reg  signReg_249; // @[block_division.scala 205:28]
  wire [9:0] multiplication_249 = multiplierReg_249 * io_man_b_249; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_57_T_23 = multiplication_249 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_249; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_57_T_22 = {1'h0,dotProductRegs_3_57}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_57_T_23 = ~_two_complement_57_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_57_T_25 = _two_complement_57_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_250; // @[block_division.scala 204:34]
  reg  signReg_250; // @[block_division.scala 205:28]
  wire [9:0] multiplication_250 = multiplierReg_250 * io_man_b_250; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_58_T_23 = multiplication_250 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_250; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_58_T_22 = {1'h0,dotProductRegs_3_58}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_58_T_23 = ~_two_complement_58_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_58_T_25 = _two_complement_58_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_251; // @[block_division.scala 204:34]
  reg  signReg_251; // @[block_division.scala 205:28]
  wire [9:0] multiplication_251 = multiplierReg_251 * io_man_b_251; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_59_T_23 = multiplication_251 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_251; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_59_T_22 = {1'h0,dotProductRegs_3_59}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_59_T_23 = ~_two_complement_59_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_59_T_25 = _two_complement_59_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_252; // @[block_division.scala 204:34]
  reg  signReg_252; // @[block_division.scala 205:28]
  wire [9:0] multiplication_252 = multiplierReg_252 * io_man_b_252; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_60_T_23 = multiplication_252 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_252; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_60_T_22 = {1'h0,dotProductRegs_3_60}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_60_T_23 = ~_two_complement_60_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_60_T_25 = _two_complement_60_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_253; // @[block_division.scala 204:34]
  reg  signReg_253; // @[block_division.scala 205:28]
  wire [9:0] multiplication_253 = multiplierReg_253 * io_man_b_253; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_61_T_23 = multiplication_253 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_253; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_61_T_22 = {1'h0,dotProductRegs_3_61}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_61_T_23 = ~_two_complement_61_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_61_T_25 = _two_complement_61_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_254; // @[block_division.scala 204:34]
  reg  signReg_254; // @[block_division.scala 205:28]
  wire [9:0] multiplication_254 = multiplierReg_254 * io_man_b_254; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_62_T_23 = multiplication_254 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_254; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_62_T_22 = {1'h0,dotProductRegs_3_62}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_62_T_23 = ~_two_complement_62_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_62_T_25 = _two_complement_62_T_23 + 6'h1; // @[block_division.scala 213:38]
  reg [4:0] multiplierReg_255; // @[block_division.scala 204:34]
  reg  signReg_255; // @[block_division.scala 205:28]
  wire [9:0] multiplication_255 = multiplierReg_255 * io_man_b_255; // @[block_division.scala 208:42]
  wire [9:0] _dotProductRegs_63_T_23 = multiplication_255 > _GEN_0 ? {{4'd0}, _dotProductRegs_0_T_1} :
    multiplication_255; // @[block_division.scala 209:31]
  wire [5:0] _two_complement_63_T_22 = {1'h0,dotProductRegs_3_63}; // @[block_division.scala 213:16]
  wire [5:0] _two_complement_63_T_23 = ~_two_complement_63_T_22; // @[block_division.scala 213:10]
  wire [5:0] _two_complement_63_T_25 = _two_complement_63_T_23 + 6'h1; // @[block_division.scala 213:38]
  wire [6:0] _sum_T_186 = $signed(two_complement_buffer_3_0) + $signed(two_complement_buffer_3_1); // @[block_division.scala 218:46]
  wire [6:0] _GEN_448 = {{1{two_complement_buffer_3_2[5]}},two_complement_buffer_3_2}; // @[block_division.scala 218:46]
  wire [7:0] _sum_T_187 = $signed(_sum_T_186) + $signed(_GEN_448); // @[block_division.scala 218:46]
  wire [7:0] _GEN_449 = {{2{two_complement_buffer_3_3[5]}},two_complement_buffer_3_3}; // @[block_division.scala 218:46]
  wire [8:0] _sum_T_188 = $signed(_sum_T_187) + $signed(_GEN_449); // @[block_division.scala 218:46]
  wire [8:0] _GEN_450 = {{3{two_complement_buffer_3_4[5]}},two_complement_buffer_3_4}; // @[block_division.scala 218:46]
  wire [9:0] _sum_T_189 = $signed(_sum_T_188) + $signed(_GEN_450); // @[block_division.scala 218:46]
  wire [9:0] _GEN_451 = {{4{two_complement_buffer_3_5[5]}},two_complement_buffer_3_5}; // @[block_division.scala 218:46]
  wire [10:0] _sum_T_190 = $signed(_sum_T_189) + $signed(_GEN_451); // @[block_division.scala 218:46]
  wire [10:0] _GEN_452 = {{5{two_complement_buffer_3_6[5]}},two_complement_buffer_3_6}; // @[block_division.scala 218:46]
  wire [11:0] _sum_T_191 = $signed(_sum_T_190) + $signed(_GEN_452); // @[block_division.scala 218:46]
  wire [11:0] _GEN_453 = {{6{two_complement_buffer_3_7[5]}},two_complement_buffer_3_7}; // @[block_division.scala 218:46]
  wire [12:0] _sum_T_192 = $signed(_sum_T_191) + $signed(_GEN_453); // @[block_division.scala 218:46]
  wire [12:0] _GEN_454 = {{7{two_complement_buffer_3_8[5]}},two_complement_buffer_3_8}; // @[block_division.scala 218:46]
  wire [13:0] _sum_T_193 = $signed(_sum_T_192) + $signed(_GEN_454); // @[block_division.scala 218:46]
  wire [13:0] _GEN_455 = {{8{two_complement_buffer_3_9[5]}},two_complement_buffer_3_9}; // @[block_division.scala 218:46]
  wire [14:0] _sum_T_194 = $signed(_sum_T_193) + $signed(_GEN_455); // @[block_division.scala 218:46]
  wire [14:0] _GEN_456 = {{9{two_complement_buffer_3_10[5]}},two_complement_buffer_3_10}; // @[block_division.scala 218:46]
  wire [15:0] _sum_T_195 = $signed(_sum_T_194) + $signed(_GEN_456); // @[block_division.scala 218:46]
  wire [15:0] _GEN_457 = {{10{two_complement_buffer_3_11[5]}},two_complement_buffer_3_11}; // @[block_division.scala 218:46]
  wire [16:0] _sum_T_196 = $signed(_sum_T_195) + $signed(_GEN_457); // @[block_division.scala 218:46]
  wire [16:0] _GEN_458 = {{11{two_complement_buffer_3_12[5]}},two_complement_buffer_3_12}; // @[block_division.scala 218:46]
  wire [17:0] _sum_T_197 = $signed(_sum_T_196) + $signed(_GEN_458); // @[block_division.scala 218:46]
  wire [17:0] _GEN_459 = {{12{two_complement_buffer_3_13[5]}},two_complement_buffer_3_13}; // @[block_division.scala 218:46]
  wire [18:0] _sum_T_198 = $signed(_sum_T_197) + $signed(_GEN_459); // @[block_division.scala 218:46]
  wire [18:0] _GEN_460 = {{13{two_complement_buffer_3_14[5]}},two_complement_buffer_3_14}; // @[block_division.scala 218:46]
  wire [19:0] _sum_T_199 = $signed(_sum_T_198) + $signed(_GEN_460); // @[block_division.scala 218:46]
  wire [19:0] _GEN_461 = {{14{two_complement_buffer_3_15[5]}},two_complement_buffer_3_15}; // @[block_division.scala 218:46]
  wire [20:0] _sum_T_200 = $signed(_sum_T_199) + $signed(_GEN_461); // @[block_division.scala 218:46]
  wire [20:0] _GEN_462 = {{15{two_complement_buffer_3_16[5]}},two_complement_buffer_3_16}; // @[block_division.scala 218:46]
  wire [21:0] _sum_T_201 = $signed(_sum_T_200) + $signed(_GEN_462); // @[block_division.scala 218:46]
  wire [21:0] _GEN_463 = {{16{two_complement_buffer_3_17[5]}},two_complement_buffer_3_17}; // @[block_division.scala 218:46]
  wire [22:0] _sum_T_202 = $signed(_sum_T_201) + $signed(_GEN_463); // @[block_division.scala 218:46]
  wire [22:0] _GEN_464 = {{17{two_complement_buffer_3_18[5]}},two_complement_buffer_3_18}; // @[block_division.scala 218:46]
  wire [23:0] _sum_T_203 = $signed(_sum_T_202) + $signed(_GEN_464); // @[block_division.scala 218:46]
  wire [23:0] _GEN_465 = {{18{two_complement_buffer_3_19[5]}},two_complement_buffer_3_19}; // @[block_division.scala 218:46]
  wire [24:0] _sum_T_204 = $signed(_sum_T_203) + $signed(_GEN_465); // @[block_division.scala 218:46]
  wire [24:0] _GEN_466 = {{19{two_complement_buffer_3_20[5]}},two_complement_buffer_3_20}; // @[block_division.scala 218:46]
  wire [25:0] _sum_T_205 = $signed(_sum_T_204) + $signed(_GEN_466); // @[block_division.scala 218:46]
  wire [25:0] _GEN_467 = {{20{two_complement_buffer_3_21[5]}},two_complement_buffer_3_21}; // @[block_division.scala 218:46]
  wire [26:0] _sum_T_206 = $signed(_sum_T_205) + $signed(_GEN_467); // @[block_division.scala 218:46]
  wire [26:0] _GEN_468 = {{21{two_complement_buffer_3_22[5]}},two_complement_buffer_3_22}; // @[block_division.scala 218:46]
  wire [27:0] _sum_T_207 = $signed(_sum_T_206) + $signed(_GEN_468); // @[block_division.scala 218:46]
  wire [27:0] _GEN_469 = {{22{two_complement_buffer_3_23[5]}},two_complement_buffer_3_23}; // @[block_division.scala 218:46]
  wire [28:0] _sum_T_208 = $signed(_sum_T_207) + $signed(_GEN_469); // @[block_division.scala 218:46]
  wire [28:0] _GEN_470 = {{23{two_complement_buffer_3_24[5]}},two_complement_buffer_3_24}; // @[block_division.scala 218:46]
  wire [29:0] _sum_T_209 = $signed(_sum_T_208) + $signed(_GEN_470); // @[block_division.scala 218:46]
  wire [29:0] _GEN_471 = {{24{two_complement_buffer_3_25[5]}},two_complement_buffer_3_25}; // @[block_division.scala 218:46]
  wire [30:0] _sum_T_210 = $signed(_sum_T_209) + $signed(_GEN_471); // @[block_division.scala 218:46]
  wire [30:0] _GEN_472 = {{25{two_complement_buffer_3_26[5]}},two_complement_buffer_3_26}; // @[block_division.scala 218:46]
  wire [31:0] _sum_T_211 = $signed(_sum_T_210) + $signed(_GEN_472); // @[block_division.scala 218:46]
  wire [31:0] _GEN_473 = {{26{two_complement_buffer_3_27[5]}},two_complement_buffer_3_27}; // @[block_division.scala 218:46]
  wire [32:0] _sum_T_212 = $signed(_sum_T_211) + $signed(_GEN_473); // @[block_division.scala 218:46]
  wire [32:0] _GEN_474 = {{27{two_complement_buffer_3_28[5]}},two_complement_buffer_3_28}; // @[block_division.scala 218:46]
  wire [33:0] _sum_T_213 = $signed(_sum_T_212) + $signed(_GEN_474); // @[block_division.scala 218:46]
  wire [33:0] _GEN_475 = {{28{two_complement_buffer_3_29[5]}},two_complement_buffer_3_29}; // @[block_division.scala 218:46]
  wire [34:0] _sum_T_214 = $signed(_sum_T_213) + $signed(_GEN_475); // @[block_division.scala 218:46]
  wire [34:0] _GEN_476 = {{29{two_complement_buffer_3_30[5]}},two_complement_buffer_3_30}; // @[block_division.scala 218:46]
  wire [35:0] _sum_T_215 = $signed(_sum_T_214) + $signed(_GEN_476); // @[block_division.scala 218:46]
  wire [35:0] _GEN_477 = {{30{two_complement_buffer_3_31[5]}},two_complement_buffer_3_31}; // @[block_division.scala 218:46]
  wire [36:0] _sum_T_216 = $signed(_sum_T_215) + $signed(_GEN_477); // @[block_division.scala 218:46]
  wire [36:0] _GEN_478 = {{31{two_complement_buffer_3_32[5]}},two_complement_buffer_3_32}; // @[block_division.scala 218:46]
  wire [37:0] _sum_T_217 = $signed(_sum_T_216) + $signed(_GEN_478); // @[block_division.scala 218:46]
  wire [37:0] _GEN_479 = {{32{two_complement_buffer_3_33[5]}},two_complement_buffer_3_33}; // @[block_division.scala 218:46]
  wire [38:0] _sum_T_218 = $signed(_sum_T_217) + $signed(_GEN_479); // @[block_division.scala 218:46]
  wire [38:0] _GEN_480 = {{33{two_complement_buffer_3_34[5]}},two_complement_buffer_3_34}; // @[block_division.scala 218:46]
  wire [39:0] _sum_T_219 = $signed(_sum_T_218) + $signed(_GEN_480); // @[block_division.scala 218:46]
  wire [39:0] _GEN_481 = {{34{two_complement_buffer_3_35[5]}},two_complement_buffer_3_35}; // @[block_division.scala 218:46]
  wire [40:0] _sum_T_220 = $signed(_sum_T_219) + $signed(_GEN_481); // @[block_division.scala 218:46]
  wire [40:0] _GEN_482 = {{35{two_complement_buffer_3_36[5]}},two_complement_buffer_3_36}; // @[block_division.scala 218:46]
  wire [41:0] _sum_T_221 = $signed(_sum_T_220) + $signed(_GEN_482); // @[block_division.scala 218:46]
  wire [41:0] _GEN_483 = {{36{two_complement_buffer_3_37[5]}},two_complement_buffer_3_37}; // @[block_division.scala 218:46]
  wire [42:0] _sum_T_222 = $signed(_sum_T_221) + $signed(_GEN_483); // @[block_division.scala 218:46]
  wire [42:0] _GEN_484 = {{37{two_complement_buffer_3_38[5]}},two_complement_buffer_3_38}; // @[block_division.scala 218:46]
  wire [43:0] _sum_T_223 = $signed(_sum_T_222) + $signed(_GEN_484); // @[block_division.scala 218:46]
  wire [43:0] _GEN_485 = {{38{two_complement_buffer_3_39[5]}},two_complement_buffer_3_39}; // @[block_division.scala 218:46]
  wire [44:0] _sum_T_224 = $signed(_sum_T_223) + $signed(_GEN_485); // @[block_division.scala 218:46]
  wire [44:0] _GEN_486 = {{39{two_complement_buffer_3_40[5]}},two_complement_buffer_3_40}; // @[block_division.scala 218:46]
  wire [45:0] _sum_T_225 = $signed(_sum_T_224) + $signed(_GEN_486); // @[block_division.scala 218:46]
  wire [45:0] _GEN_487 = {{40{two_complement_buffer_3_41[5]}},two_complement_buffer_3_41}; // @[block_division.scala 218:46]
  wire [46:0] _sum_T_226 = $signed(_sum_T_225) + $signed(_GEN_487); // @[block_division.scala 218:46]
  wire [46:0] _GEN_488 = {{41{two_complement_buffer_3_42[5]}},two_complement_buffer_3_42}; // @[block_division.scala 218:46]
  wire [47:0] _sum_T_227 = $signed(_sum_T_226) + $signed(_GEN_488); // @[block_division.scala 218:46]
  wire [47:0] _GEN_489 = {{42{two_complement_buffer_3_43[5]}},two_complement_buffer_3_43}; // @[block_division.scala 218:46]
  wire [48:0] _sum_T_228 = $signed(_sum_T_227) + $signed(_GEN_489); // @[block_division.scala 218:46]
  wire [48:0] _GEN_490 = {{43{two_complement_buffer_3_44[5]}},two_complement_buffer_3_44}; // @[block_division.scala 218:46]
  wire [49:0] _sum_T_229 = $signed(_sum_T_228) + $signed(_GEN_490); // @[block_division.scala 218:46]
  wire [49:0] _GEN_491 = {{44{two_complement_buffer_3_45[5]}},two_complement_buffer_3_45}; // @[block_division.scala 218:46]
  wire [50:0] _sum_T_230 = $signed(_sum_T_229) + $signed(_GEN_491); // @[block_division.scala 218:46]
  wire [50:0] _GEN_492 = {{45{two_complement_buffer_3_46[5]}},two_complement_buffer_3_46}; // @[block_division.scala 218:46]
  wire [51:0] _sum_T_231 = $signed(_sum_T_230) + $signed(_GEN_492); // @[block_division.scala 218:46]
  wire [51:0] _GEN_493 = {{46{two_complement_buffer_3_47[5]}},two_complement_buffer_3_47}; // @[block_division.scala 218:46]
  wire [52:0] _sum_T_232 = $signed(_sum_T_231) + $signed(_GEN_493); // @[block_division.scala 218:46]
  wire [52:0] _GEN_494 = {{47{two_complement_buffer_3_48[5]}},two_complement_buffer_3_48}; // @[block_division.scala 218:46]
  wire [53:0] _sum_T_233 = $signed(_sum_T_232) + $signed(_GEN_494); // @[block_division.scala 218:46]
  wire [53:0] _GEN_495 = {{48{two_complement_buffer_3_49[5]}},two_complement_buffer_3_49}; // @[block_division.scala 218:46]
  wire [54:0] _sum_T_234 = $signed(_sum_T_233) + $signed(_GEN_495); // @[block_division.scala 218:46]
  wire [54:0] _GEN_496 = {{49{two_complement_buffer_3_50[5]}},two_complement_buffer_3_50}; // @[block_division.scala 218:46]
  wire [55:0] _sum_T_235 = $signed(_sum_T_234) + $signed(_GEN_496); // @[block_division.scala 218:46]
  wire [55:0] _GEN_497 = {{50{two_complement_buffer_3_51[5]}},two_complement_buffer_3_51}; // @[block_division.scala 218:46]
  wire [56:0] _sum_T_236 = $signed(_sum_T_235) + $signed(_GEN_497); // @[block_division.scala 218:46]
  wire [56:0] _GEN_498 = {{51{two_complement_buffer_3_52[5]}},two_complement_buffer_3_52}; // @[block_division.scala 218:46]
  wire [57:0] _sum_T_237 = $signed(_sum_T_236) + $signed(_GEN_498); // @[block_division.scala 218:46]
  wire [57:0] _GEN_499 = {{52{two_complement_buffer_3_53[5]}},two_complement_buffer_3_53}; // @[block_division.scala 218:46]
  wire [58:0] _sum_T_238 = $signed(_sum_T_237) + $signed(_GEN_499); // @[block_division.scala 218:46]
  wire [58:0] _GEN_500 = {{53{two_complement_buffer_3_54[5]}},two_complement_buffer_3_54}; // @[block_division.scala 218:46]
  wire [59:0] _sum_T_239 = $signed(_sum_T_238) + $signed(_GEN_500); // @[block_division.scala 218:46]
  wire [59:0] _GEN_501 = {{54{two_complement_buffer_3_55[5]}},two_complement_buffer_3_55}; // @[block_division.scala 218:46]
  wire [60:0] _sum_T_240 = $signed(_sum_T_239) + $signed(_GEN_501); // @[block_division.scala 218:46]
  wire [60:0] _GEN_502 = {{55{two_complement_buffer_3_56[5]}},two_complement_buffer_3_56}; // @[block_division.scala 218:46]
  wire [61:0] _sum_T_241 = $signed(_sum_T_240) + $signed(_GEN_502); // @[block_division.scala 218:46]
  wire [61:0] _GEN_503 = {{56{two_complement_buffer_3_57[5]}},two_complement_buffer_3_57}; // @[block_division.scala 218:46]
  wire [62:0] _sum_T_242 = $signed(_sum_T_241) + $signed(_GEN_503); // @[block_division.scala 218:46]
  wire [62:0] _GEN_504 = {{57{two_complement_buffer_3_58[5]}},two_complement_buffer_3_58}; // @[block_division.scala 218:46]
  wire [63:0] _sum_T_243 = $signed(_sum_T_242) + $signed(_GEN_504); // @[block_division.scala 218:46]
  wire [63:0] _GEN_505 = {{58{two_complement_buffer_3_59[5]}},two_complement_buffer_3_59}; // @[block_division.scala 218:46]
  wire [64:0] _sum_T_244 = $signed(_sum_T_243) + $signed(_GEN_505); // @[block_division.scala 218:46]
  wire [64:0] _GEN_506 = {{59{two_complement_buffer_3_60[5]}},two_complement_buffer_3_60}; // @[block_division.scala 218:46]
  wire [65:0] _sum_T_245 = $signed(_sum_T_244) + $signed(_GEN_506); // @[block_division.scala 218:46]
  wire [65:0] _GEN_507 = {{60{two_complement_buffer_3_61[5]}},two_complement_buffer_3_61}; // @[block_division.scala 218:46]
  wire [66:0] _sum_T_246 = $signed(_sum_T_245) + $signed(_GEN_507); // @[block_division.scala 218:46]
  wire [66:0] _GEN_508 = {{61{two_complement_buffer_3_62[5]}},two_complement_buffer_3_62}; // @[block_division.scala 218:46]
  wire [67:0] _sum_T_247 = $signed(_sum_T_246) + $signed(_GEN_508); // @[block_division.scala 218:46]
  wire [67:0] _GEN_509 = {{62{two_complement_buffer_3_63[5]}},two_complement_buffer_3_63}; // @[block_division.scala 218:46]
  wire [68:0] sum_3 = $signed(_sum_T_247) + $signed(_GEN_509); // @[block_division.scala 218:46]
  wire [67:0] _acc_3_T_3 = ~sum_3[67:0]; // @[block_division.scala 219:57]
  wire [67:0] _acc_3_T_5 = _acc_3_T_3 + 68'h1; // @[block_division.scala 219:86]
  wire [68:0] _acc_3_T_14 = $signed(_sum_T_247) + $signed(_GEN_509); // @[block_division.scala 219:145]
  wire [68:0] _acc_3_T_15 = _acc_3_T_5 > _GEN_126 ? {{63'd0}, _acc_0_T_13} : _acc_3_T_14; // @[block_division.scala 219:55]
  wire [68:0] _acc_3_T_23 = sum_3[67:0] > _GEN_126 ? {{63'd0}, _dotProductRegs_0_T_1} : _acc_3_T_14; // @[block_division.scala 220:6]
  wire [68:0] _acc_3_T_24 = sum_3[68] ? _acc_3_T_15 : _acc_3_T_23; // @[block_division.scala 219:18]
  wire [68:0] _GEN_512 = reset ? 69'h0 : _acc_0_T_24; // @[block_division.scala 195:{53,53} 219:12]
  wire [68:0] _GEN_513 = reset ? 69'h0 : _acc_1_T_24; // @[block_division.scala 195:{53,53} 219:12]
  wire [68:0] _GEN_514 = reset ? 69'h0 : _acc_2_T_24; // @[block_division.scala 195:{53,53} 219:12]
  wire [68:0] _GEN_515 = reset ? 69'h0 : _acc_3_T_24; // @[block_division.scala 195:{53,53} 219:12]
  adderTree2 adderTreeInst ( // @[block_division.scala 223:29]
    .clock(adderTreeInst_clock),
    .reset(adderTreeInst_reset),
    .io_sign_man_0(adderTreeInst_io_sign_man_0),
    .io_sign_man_1(adderTreeInst_io_sign_man_1),
    .io_sign_man_2(adderTreeInst_io_sign_man_2),
    .io_sign_man_3(adderTreeInst_io_sign_man_3),
    .io_exps_0(adderTreeInst_io_exps_0),
    .io_exps_1(adderTreeInst_io_exps_1),
    .io_exps_2(adderTreeInst_io_exps_2),
    .io_exps_3(adderTreeInst_io_exps_3),
    .io_control_signal(adderTreeInst_io_control_signal),
    .io_control_signal2(adderTreeInst_io_control_signal2),
    .io_result_tree(adderTreeInst_io_result_tree)
  );
  assign io_result = adderTreeInst_io_result_tree; // @[block_division.scala 228:13]
  assign adderTreeInst_clock = clock;
  assign adderTreeInst_reset = reset;
  assign adderTreeInst_io_sign_man_0 = acc_0; // @[block_division.scala 224:{39,39}]
  assign adderTreeInst_io_sign_man_1 = acc_1; // @[block_division.scala 224:{39,39}]
  assign adderTreeInst_io_sign_man_2 = acc_2; // @[block_division.scala 224:{39,39}]
  assign adderTreeInst_io_sign_man_3 = acc_3; // @[block_division.scala 224:{39,39}]
  assign adderTreeInst_io_exps_0 = exp_output_0; // @[block_division.scala 225:{35,35}]
  assign adderTreeInst_io_exps_1 = exp_output_1; // @[block_division.scala 225:{35,35}]
  assign adderTreeInst_io_exps_2 = exp_output_2; // @[block_division.scala 225:{35,35}]
  assign adderTreeInst_io_exps_3 = exp_output_3; // @[block_division.scala 225:{35,35}]
  assign adderTreeInst_io_control_signal = io_control; // @[block_division.scala 226:35]
  assign adderTreeInst_io_control_signal2 = io_control2; // @[block_division.scala 227:36]
  always @(posedge clock) begin
    if (reset) begin // @[block_division.scala 194:60]
      exp_output_0 <= 9'h0; // @[block_division.scala 194:60]
    end else begin
      exp_output_0 <= _exp_output_0_T; // @[block_division.scala 198:19]
    end
    if (reset) begin // @[block_division.scala 194:60]
      exp_output_1 <= 9'h0; // @[block_division.scala 194:60]
    end else begin
      exp_output_1 <= _exp_output_1_T; // @[block_division.scala 198:19]
    end
    if (reset) begin // @[block_division.scala 194:60]
      exp_output_2 <= 9'h0; // @[block_division.scala 194:60]
    end else begin
      exp_output_2 <= _exp_output_2_T; // @[block_division.scala 198:19]
    end
    if (reset) begin // @[block_division.scala 194:60]
      exp_output_3 <= 9'h0; // @[block_division.scala 194:60]
    end else begin
      exp_output_3 <= _exp_output_3_T; // @[block_division.scala 198:19]
    end
    acc_0 <= _GEN_512[5:0]; // @[block_division.scala 195:{53,53} 219:12]
    acc_1 <= _GEN_513[5:0]; // @[block_division.scala 195:{53,53} 219:12]
    acc_2 <= _GEN_514[5:0]; // @[block_division.scala 195:{53,53} 219:12]
    acc_3 <= _GEN_515[5:0]; // @[block_division.scala 195:{53,53} 219:12]
    dotProductRegs__0 <= _dotProductRegs_0_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__1 <= _dotProductRegs_1_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__2 <= _dotProductRegs_2_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__3 <= _dotProductRegs_3_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__4 <= _dotProductRegs_4_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__5 <= _dotProductRegs_5_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__6 <= _dotProductRegs_6_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__7 <= _dotProductRegs_7_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__8 <= _dotProductRegs_8_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__9 <= _dotProductRegs_9_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__10 <= _dotProductRegs_10_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__11 <= _dotProductRegs_11_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__12 <= _dotProductRegs_12_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__13 <= _dotProductRegs_13_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__14 <= _dotProductRegs_14_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__15 <= _dotProductRegs_15_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__16 <= _dotProductRegs_16_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__17 <= _dotProductRegs_17_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__18 <= _dotProductRegs_18_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__19 <= _dotProductRegs_19_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__20 <= _dotProductRegs_20_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__21 <= _dotProductRegs_21_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__22 <= _dotProductRegs_22_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__23 <= _dotProductRegs_23_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__24 <= _dotProductRegs_24_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__25 <= _dotProductRegs_25_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__26 <= _dotProductRegs_26_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__27 <= _dotProductRegs_27_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__28 <= _dotProductRegs_28_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__29 <= _dotProductRegs_29_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__30 <= _dotProductRegs_30_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__31 <= _dotProductRegs_31_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__32 <= _dotProductRegs_32_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__33 <= _dotProductRegs_33_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__34 <= _dotProductRegs_34_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__35 <= _dotProductRegs_35_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__36 <= _dotProductRegs_36_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__37 <= _dotProductRegs_37_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__38 <= _dotProductRegs_38_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__39 <= _dotProductRegs_39_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__40 <= _dotProductRegs_40_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__41 <= _dotProductRegs_41_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__42 <= _dotProductRegs_42_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__43 <= _dotProductRegs_43_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__44 <= _dotProductRegs_44_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__45 <= _dotProductRegs_45_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__46 <= _dotProductRegs_46_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__47 <= _dotProductRegs_47_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__48 <= _dotProductRegs_48_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__49 <= _dotProductRegs_49_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__50 <= _dotProductRegs_50_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__51 <= _dotProductRegs_51_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__52 <= _dotProductRegs_52_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__53 <= _dotProductRegs_53_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__54 <= _dotProductRegs_54_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__55 <= _dotProductRegs_55_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__56 <= _dotProductRegs_56_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__57 <= _dotProductRegs_57_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__58 <= _dotProductRegs_58_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__59 <= _dotProductRegs_59_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__60 <= _dotProductRegs_60_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__61 <= _dotProductRegs_61_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__62 <= _dotProductRegs_62_T_5[4:0]; // @[block_division.scala 209:25]
    dotProductRegs__63 <= _dotProductRegs_63_T_5[4:0]; // @[block_division.scala 209:25]
    signs__0 <= signReg ^ io_sign_b_0; // @[block_division.scala 210:27]
    signs__1 <= signReg_1 ^ io_sign_b_1; // @[block_division.scala 210:27]
    signs__2 <= signReg_2 ^ io_sign_b_2; // @[block_division.scala 210:27]
    signs__3 <= signReg_3 ^ io_sign_b_3; // @[block_division.scala 210:27]
    signs__4 <= signReg_4 ^ io_sign_b_4; // @[block_division.scala 210:27]
    signs__5 <= signReg_5 ^ io_sign_b_5; // @[block_division.scala 210:27]
    signs__6 <= signReg_6 ^ io_sign_b_6; // @[block_division.scala 210:27]
    signs__7 <= signReg_7 ^ io_sign_b_7; // @[block_division.scala 210:27]
    signs__8 <= signReg_8 ^ io_sign_b_8; // @[block_division.scala 210:27]
    signs__9 <= signReg_9 ^ io_sign_b_9; // @[block_division.scala 210:27]
    signs__10 <= signReg_10 ^ io_sign_b_10; // @[block_division.scala 210:27]
    signs__11 <= signReg_11 ^ io_sign_b_11; // @[block_division.scala 210:27]
    signs__12 <= signReg_12 ^ io_sign_b_12; // @[block_division.scala 210:27]
    signs__13 <= signReg_13 ^ io_sign_b_13; // @[block_division.scala 210:27]
    signs__14 <= signReg_14 ^ io_sign_b_14; // @[block_division.scala 210:27]
    signs__15 <= signReg_15 ^ io_sign_b_15; // @[block_division.scala 210:27]
    signs__16 <= signReg_16 ^ io_sign_b_16; // @[block_division.scala 210:27]
    signs__17 <= signReg_17 ^ io_sign_b_17; // @[block_division.scala 210:27]
    signs__18 <= signReg_18 ^ io_sign_b_18; // @[block_division.scala 210:27]
    signs__19 <= signReg_19 ^ io_sign_b_19; // @[block_division.scala 210:27]
    signs__20 <= signReg_20 ^ io_sign_b_20; // @[block_division.scala 210:27]
    signs__21 <= signReg_21 ^ io_sign_b_21; // @[block_division.scala 210:27]
    signs__22 <= signReg_22 ^ io_sign_b_22; // @[block_division.scala 210:27]
    signs__23 <= signReg_23 ^ io_sign_b_23; // @[block_division.scala 210:27]
    signs__24 <= signReg_24 ^ io_sign_b_24; // @[block_division.scala 210:27]
    signs__25 <= signReg_25 ^ io_sign_b_25; // @[block_division.scala 210:27]
    signs__26 <= signReg_26 ^ io_sign_b_26; // @[block_division.scala 210:27]
    signs__27 <= signReg_27 ^ io_sign_b_27; // @[block_division.scala 210:27]
    signs__28 <= signReg_28 ^ io_sign_b_28; // @[block_division.scala 210:27]
    signs__29 <= signReg_29 ^ io_sign_b_29; // @[block_division.scala 210:27]
    signs__30 <= signReg_30 ^ io_sign_b_30; // @[block_division.scala 210:27]
    signs__31 <= signReg_31 ^ io_sign_b_31; // @[block_division.scala 210:27]
    signs__32 <= signReg_32 ^ io_sign_b_32; // @[block_division.scala 210:27]
    signs__33 <= signReg_33 ^ io_sign_b_33; // @[block_division.scala 210:27]
    signs__34 <= signReg_34 ^ io_sign_b_34; // @[block_division.scala 210:27]
    signs__35 <= signReg_35 ^ io_sign_b_35; // @[block_division.scala 210:27]
    signs__36 <= signReg_36 ^ io_sign_b_36; // @[block_division.scala 210:27]
    signs__37 <= signReg_37 ^ io_sign_b_37; // @[block_division.scala 210:27]
    signs__38 <= signReg_38 ^ io_sign_b_38; // @[block_division.scala 210:27]
    signs__39 <= signReg_39 ^ io_sign_b_39; // @[block_division.scala 210:27]
    signs__40 <= signReg_40 ^ io_sign_b_40; // @[block_division.scala 210:27]
    signs__41 <= signReg_41 ^ io_sign_b_41; // @[block_division.scala 210:27]
    signs__42 <= signReg_42 ^ io_sign_b_42; // @[block_division.scala 210:27]
    signs__43 <= signReg_43 ^ io_sign_b_43; // @[block_division.scala 210:27]
    signs__44 <= signReg_44 ^ io_sign_b_44; // @[block_division.scala 210:27]
    signs__45 <= signReg_45 ^ io_sign_b_45; // @[block_division.scala 210:27]
    signs__46 <= signReg_46 ^ io_sign_b_46; // @[block_division.scala 210:27]
    signs__47 <= signReg_47 ^ io_sign_b_47; // @[block_division.scala 210:27]
    signs__48 <= signReg_48 ^ io_sign_b_48; // @[block_division.scala 210:27]
    signs__49 <= signReg_49 ^ io_sign_b_49; // @[block_division.scala 210:27]
    signs__50 <= signReg_50 ^ io_sign_b_50; // @[block_division.scala 210:27]
    signs__51 <= signReg_51 ^ io_sign_b_51; // @[block_division.scala 210:27]
    signs__52 <= signReg_52 ^ io_sign_b_52; // @[block_division.scala 210:27]
    signs__53 <= signReg_53 ^ io_sign_b_53; // @[block_division.scala 210:27]
    signs__54 <= signReg_54 ^ io_sign_b_54; // @[block_division.scala 210:27]
    signs__55 <= signReg_55 ^ io_sign_b_55; // @[block_division.scala 210:27]
    signs__56 <= signReg_56 ^ io_sign_b_56; // @[block_division.scala 210:27]
    signs__57 <= signReg_57 ^ io_sign_b_57; // @[block_division.scala 210:27]
    signs__58 <= signReg_58 ^ io_sign_b_58; // @[block_division.scala 210:27]
    signs__59 <= signReg_59 ^ io_sign_b_59; // @[block_division.scala 210:27]
    signs__60 <= signReg_60 ^ io_sign_b_60; // @[block_division.scala 210:27]
    signs__61 <= signReg_61 ^ io_sign_b_61; // @[block_division.scala 210:27]
    signs__62 <= signReg_62 ^ io_sign_b_62; // @[block_division.scala 210:27]
    signs__63 <= signReg_63 ^ io_sign_b_63; // @[block_division.scala 210:27]
    if (signs__0) begin // @[block_division.scala 211:31]
      two_complement__0 <= _two_complement_0_T_4;
    end else begin
      two_complement__0 <= _two_complement_0_T_1;
    end
    if (signs__1) begin // @[block_division.scala 211:31]
      two_complement__1 <= _two_complement_1_T_4;
    end else begin
      two_complement__1 <= _two_complement_1_T_1;
    end
    if (signs__2) begin // @[block_division.scala 211:31]
      two_complement__2 <= _two_complement_2_T_4;
    end else begin
      two_complement__2 <= _two_complement_2_T_1;
    end
    if (signs__3) begin // @[block_division.scala 211:31]
      two_complement__3 <= _two_complement_3_T_4;
    end else begin
      two_complement__3 <= _two_complement_3_T_1;
    end
    if (signs__4) begin // @[block_division.scala 211:31]
      two_complement__4 <= _two_complement_4_T_4;
    end else begin
      two_complement__4 <= _two_complement_4_T_1;
    end
    if (signs__5) begin // @[block_division.scala 211:31]
      two_complement__5 <= _two_complement_5_T_4;
    end else begin
      two_complement__5 <= _two_complement_5_T_1;
    end
    if (signs__6) begin // @[block_division.scala 211:31]
      two_complement__6 <= _two_complement_6_T_4;
    end else begin
      two_complement__6 <= _two_complement_6_T_1;
    end
    if (signs__7) begin // @[block_division.scala 211:31]
      two_complement__7 <= _two_complement_7_T_4;
    end else begin
      two_complement__7 <= _two_complement_7_T_1;
    end
    if (signs__8) begin // @[block_division.scala 211:31]
      two_complement__8 <= _two_complement_8_T_4;
    end else begin
      two_complement__8 <= _two_complement_8_T_1;
    end
    if (signs__9) begin // @[block_division.scala 211:31]
      two_complement__9 <= _two_complement_9_T_4;
    end else begin
      two_complement__9 <= _two_complement_9_T_1;
    end
    if (signs__10) begin // @[block_division.scala 211:31]
      two_complement__10 <= _two_complement_10_T_4;
    end else begin
      two_complement__10 <= _two_complement_10_T_1;
    end
    if (signs__11) begin // @[block_division.scala 211:31]
      two_complement__11 <= _two_complement_11_T_4;
    end else begin
      two_complement__11 <= _two_complement_11_T_1;
    end
    if (signs__12) begin // @[block_division.scala 211:31]
      two_complement__12 <= _two_complement_12_T_4;
    end else begin
      two_complement__12 <= _two_complement_12_T_1;
    end
    if (signs__13) begin // @[block_division.scala 211:31]
      two_complement__13 <= _two_complement_13_T_4;
    end else begin
      two_complement__13 <= _two_complement_13_T_1;
    end
    if (signs__14) begin // @[block_division.scala 211:31]
      two_complement__14 <= _two_complement_14_T_4;
    end else begin
      two_complement__14 <= _two_complement_14_T_1;
    end
    if (signs__15) begin // @[block_division.scala 211:31]
      two_complement__15 <= _two_complement_15_T_4;
    end else begin
      two_complement__15 <= _two_complement_15_T_1;
    end
    if (signs__16) begin // @[block_division.scala 211:31]
      two_complement__16 <= _two_complement_16_T_4;
    end else begin
      two_complement__16 <= _two_complement_16_T_1;
    end
    if (signs__17) begin // @[block_division.scala 211:31]
      two_complement__17 <= _two_complement_17_T_4;
    end else begin
      two_complement__17 <= _two_complement_17_T_1;
    end
    if (signs__18) begin // @[block_division.scala 211:31]
      two_complement__18 <= _two_complement_18_T_4;
    end else begin
      two_complement__18 <= _two_complement_18_T_1;
    end
    if (signs__19) begin // @[block_division.scala 211:31]
      two_complement__19 <= _two_complement_19_T_4;
    end else begin
      two_complement__19 <= _two_complement_19_T_1;
    end
    if (signs__20) begin // @[block_division.scala 211:31]
      two_complement__20 <= _two_complement_20_T_4;
    end else begin
      two_complement__20 <= _two_complement_20_T_1;
    end
    if (signs__21) begin // @[block_division.scala 211:31]
      two_complement__21 <= _two_complement_21_T_4;
    end else begin
      two_complement__21 <= _two_complement_21_T_1;
    end
    if (signs__22) begin // @[block_division.scala 211:31]
      two_complement__22 <= _two_complement_22_T_4;
    end else begin
      two_complement__22 <= _two_complement_22_T_1;
    end
    if (signs__23) begin // @[block_division.scala 211:31]
      two_complement__23 <= _two_complement_23_T_4;
    end else begin
      two_complement__23 <= _two_complement_23_T_1;
    end
    if (signs__24) begin // @[block_division.scala 211:31]
      two_complement__24 <= _two_complement_24_T_4;
    end else begin
      two_complement__24 <= _two_complement_24_T_1;
    end
    if (signs__25) begin // @[block_division.scala 211:31]
      two_complement__25 <= _two_complement_25_T_4;
    end else begin
      two_complement__25 <= _two_complement_25_T_1;
    end
    if (signs__26) begin // @[block_division.scala 211:31]
      two_complement__26 <= _two_complement_26_T_4;
    end else begin
      two_complement__26 <= _two_complement_26_T_1;
    end
    if (signs__27) begin // @[block_division.scala 211:31]
      two_complement__27 <= _two_complement_27_T_4;
    end else begin
      two_complement__27 <= _two_complement_27_T_1;
    end
    if (signs__28) begin // @[block_division.scala 211:31]
      two_complement__28 <= _two_complement_28_T_4;
    end else begin
      two_complement__28 <= _two_complement_28_T_1;
    end
    if (signs__29) begin // @[block_division.scala 211:31]
      two_complement__29 <= _two_complement_29_T_4;
    end else begin
      two_complement__29 <= _two_complement_29_T_1;
    end
    if (signs__30) begin // @[block_division.scala 211:31]
      two_complement__30 <= _two_complement_30_T_4;
    end else begin
      two_complement__30 <= _two_complement_30_T_1;
    end
    if (signs__31) begin // @[block_division.scala 211:31]
      two_complement__31 <= _two_complement_31_T_4;
    end else begin
      two_complement__31 <= _two_complement_31_T_1;
    end
    if (signs__32) begin // @[block_division.scala 211:31]
      two_complement__32 <= _two_complement_32_T_4;
    end else begin
      two_complement__32 <= _two_complement_32_T_1;
    end
    if (signs__33) begin // @[block_division.scala 211:31]
      two_complement__33 <= _two_complement_33_T_4;
    end else begin
      two_complement__33 <= _two_complement_33_T_1;
    end
    if (signs__34) begin // @[block_division.scala 211:31]
      two_complement__34 <= _two_complement_34_T_4;
    end else begin
      two_complement__34 <= _two_complement_34_T_1;
    end
    if (signs__35) begin // @[block_division.scala 211:31]
      two_complement__35 <= _two_complement_35_T_4;
    end else begin
      two_complement__35 <= _two_complement_35_T_1;
    end
    if (signs__36) begin // @[block_division.scala 211:31]
      two_complement__36 <= _two_complement_36_T_4;
    end else begin
      two_complement__36 <= _two_complement_36_T_1;
    end
    if (signs__37) begin // @[block_division.scala 211:31]
      two_complement__37 <= _two_complement_37_T_4;
    end else begin
      two_complement__37 <= _two_complement_37_T_1;
    end
    if (signs__38) begin // @[block_division.scala 211:31]
      two_complement__38 <= _two_complement_38_T_4;
    end else begin
      two_complement__38 <= _two_complement_38_T_1;
    end
    if (signs__39) begin // @[block_division.scala 211:31]
      two_complement__39 <= _two_complement_39_T_4;
    end else begin
      two_complement__39 <= _two_complement_39_T_1;
    end
    if (signs__40) begin // @[block_division.scala 211:31]
      two_complement__40 <= _two_complement_40_T_4;
    end else begin
      two_complement__40 <= _two_complement_40_T_1;
    end
    if (signs__41) begin // @[block_division.scala 211:31]
      two_complement__41 <= _two_complement_41_T_4;
    end else begin
      two_complement__41 <= _two_complement_41_T_1;
    end
    if (signs__42) begin // @[block_division.scala 211:31]
      two_complement__42 <= _two_complement_42_T_4;
    end else begin
      two_complement__42 <= _two_complement_42_T_1;
    end
    if (signs__43) begin // @[block_division.scala 211:31]
      two_complement__43 <= _two_complement_43_T_4;
    end else begin
      two_complement__43 <= _two_complement_43_T_1;
    end
    if (signs__44) begin // @[block_division.scala 211:31]
      two_complement__44 <= _two_complement_44_T_4;
    end else begin
      two_complement__44 <= _two_complement_44_T_1;
    end
    if (signs__45) begin // @[block_division.scala 211:31]
      two_complement__45 <= _two_complement_45_T_4;
    end else begin
      two_complement__45 <= _two_complement_45_T_1;
    end
    if (signs__46) begin // @[block_division.scala 211:31]
      two_complement__46 <= _two_complement_46_T_4;
    end else begin
      two_complement__46 <= _two_complement_46_T_1;
    end
    if (signs__47) begin // @[block_division.scala 211:31]
      two_complement__47 <= _two_complement_47_T_4;
    end else begin
      two_complement__47 <= _two_complement_47_T_1;
    end
    if (signs__48) begin // @[block_division.scala 211:31]
      two_complement__48 <= _two_complement_48_T_4;
    end else begin
      two_complement__48 <= _two_complement_48_T_1;
    end
    if (signs__49) begin // @[block_division.scala 211:31]
      two_complement__49 <= _two_complement_49_T_4;
    end else begin
      two_complement__49 <= _two_complement_49_T_1;
    end
    if (signs__50) begin // @[block_division.scala 211:31]
      two_complement__50 <= _two_complement_50_T_4;
    end else begin
      two_complement__50 <= _two_complement_50_T_1;
    end
    if (signs__51) begin // @[block_division.scala 211:31]
      two_complement__51 <= _two_complement_51_T_4;
    end else begin
      two_complement__51 <= _two_complement_51_T_1;
    end
    if (signs__52) begin // @[block_division.scala 211:31]
      two_complement__52 <= _two_complement_52_T_4;
    end else begin
      two_complement__52 <= _two_complement_52_T_1;
    end
    if (signs__53) begin // @[block_division.scala 211:31]
      two_complement__53 <= _two_complement_53_T_4;
    end else begin
      two_complement__53 <= _two_complement_53_T_1;
    end
    if (signs__54) begin // @[block_division.scala 211:31]
      two_complement__54 <= _two_complement_54_T_4;
    end else begin
      two_complement__54 <= _two_complement_54_T_1;
    end
    if (signs__55) begin // @[block_division.scala 211:31]
      two_complement__55 <= _two_complement_55_T_4;
    end else begin
      two_complement__55 <= _two_complement_55_T_1;
    end
    if (signs__56) begin // @[block_division.scala 211:31]
      two_complement__56 <= _two_complement_56_T_4;
    end else begin
      two_complement__56 <= _two_complement_56_T_1;
    end
    if (signs__57) begin // @[block_division.scala 211:31]
      two_complement__57 <= _two_complement_57_T_4;
    end else begin
      two_complement__57 <= _two_complement_57_T_1;
    end
    if (signs__58) begin // @[block_division.scala 211:31]
      two_complement__58 <= _two_complement_58_T_4;
    end else begin
      two_complement__58 <= _two_complement_58_T_1;
    end
    if (signs__59) begin // @[block_division.scala 211:31]
      two_complement__59 <= _two_complement_59_T_4;
    end else begin
      two_complement__59 <= _two_complement_59_T_1;
    end
    if (signs__60) begin // @[block_division.scala 211:31]
      two_complement__60 <= _two_complement_60_T_4;
    end else begin
      two_complement__60 <= _two_complement_60_T_1;
    end
    if (signs__61) begin // @[block_division.scala 211:31]
      two_complement__61 <= _two_complement_61_T_4;
    end else begin
      two_complement__61 <= _two_complement_61_T_1;
    end
    if (signs__62) begin // @[block_division.scala 211:31]
      two_complement__62 <= _two_complement_62_T_4;
    end else begin
      two_complement__62 <= _two_complement_62_T_1;
    end
    if (signs__63) begin // @[block_division.scala 211:31]
      two_complement__63 <= _two_complement_63_T_4;
    end else begin
      two_complement__63 <= _two_complement_63_T_1;
    end
    two_complement_buffer__0 <= two_complement__0; // @[block_division.scala 216:53]
    two_complement_buffer__1 <= two_complement__1; // @[block_division.scala 216:53]
    two_complement_buffer__2 <= two_complement__2; // @[block_division.scala 216:53]
    two_complement_buffer__3 <= two_complement__3; // @[block_division.scala 216:53]
    two_complement_buffer__4 <= two_complement__4; // @[block_division.scala 216:53]
    two_complement_buffer__5 <= two_complement__5; // @[block_division.scala 216:53]
    two_complement_buffer__6 <= two_complement__6; // @[block_division.scala 216:53]
    two_complement_buffer__7 <= two_complement__7; // @[block_division.scala 216:53]
    two_complement_buffer__8 <= two_complement__8; // @[block_division.scala 216:53]
    two_complement_buffer__9 <= two_complement__9; // @[block_division.scala 216:53]
    two_complement_buffer__10 <= two_complement__10; // @[block_division.scala 216:53]
    two_complement_buffer__11 <= two_complement__11; // @[block_division.scala 216:53]
    two_complement_buffer__12 <= two_complement__12; // @[block_division.scala 216:53]
    two_complement_buffer__13 <= two_complement__13; // @[block_division.scala 216:53]
    two_complement_buffer__14 <= two_complement__14; // @[block_division.scala 216:53]
    two_complement_buffer__15 <= two_complement__15; // @[block_division.scala 216:53]
    two_complement_buffer__16 <= two_complement__16; // @[block_division.scala 216:53]
    two_complement_buffer__17 <= two_complement__17; // @[block_division.scala 216:53]
    two_complement_buffer__18 <= two_complement__18; // @[block_division.scala 216:53]
    two_complement_buffer__19 <= two_complement__19; // @[block_division.scala 216:53]
    two_complement_buffer__20 <= two_complement__20; // @[block_division.scala 216:53]
    two_complement_buffer__21 <= two_complement__21; // @[block_division.scala 216:53]
    two_complement_buffer__22 <= two_complement__22; // @[block_division.scala 216:53]
    two_complement_buffer__23 <= two_complement__23; // @[block_division.scala 216:53]
    two_complement_buffer__24 <= two_complement__24; // @[block_division.scala 216:53]
    two_complement_buffer__25 <= two_complement__25; // @[block_division.scala 216:53]
    two_complement_buffer__26 <= two_complement__26; // @[block_division.scala 216:53]
    two_complement_buffer__27 <= two_complement__27; // @[block_division.scala 216:53]
    two_complement_buffer__28 <= two_complement__28; // @[block_division.scala 216:53]
    two_complement_buffer__29 <= two_complement__29; // @[block_division.scala 216:53]
    two_complement_buffer__30 <= two_complement__30; // @[block_division.scala 216:53]
    two_complement_buffer__31 <= two_complement__31; // @[block_division.scala 216:53]
    two_complement_buffer__32 <= two_complement__32; // @[block_division.scala 216:53]
    two_complement_buffer__33 <= two_complement__33; // @[block_division.scala 216:53]
    two_complement_buffer__34 <= two_complement__34; // @[block_division.scala 216:53]
    two_complement_buffer__35 <= two_complement__35; // @[block_division.scala 216:53]
    two_complement_buffer__36 <= two_complement__36; // @[block_division.scala 216:53]
    two_complement_buffer__37 <= two_complement__37; // @[block_division.scala 216:53]
    two_complement_buffer__38 <= two_complement__38; // @[block_division.scala 216:53]
    two_complement_buffer__39 <= two_complement__39; // @[block_division.scala 216:53]
    two_complement_buffer__40 <= two_complement__40; // @[block_division.scala 216:53]
    two_complement_buffer__41 <= two_complement__41; // @[block_division.scala 216:53]
    two_complement_buffer__42 <= two_complement__42; // @[block_division.scala 216:53]
    two_complement_buffer__43 <= two_complement__43; // @[block_division.scala 216:53]
    two_complement_buffer__44 <= two_complement__44; // @[block_division.scala 216:53]
    two_complement_buffer__45 <= two_complement__45; // @[block_division.scala 216:53]
    two_complement_buffer__46 <= two_complement__46; // @[block_division.scala 216:53]
    two_complement_buffer__47 <= two_complement__47; // @[block_division.scala 216:53]
    two_complement_buffer__48 <= two_complement__48; // @[block_division.scala 216:53]
    two_complement_buffer__49 <= two_complement__49; // @[block_division.scala 216:53]
    two_complement_buffer__50 <= two_complement__50; // @[block_division.scala 216:53]
    two_complement_buffer__51 <= two_complement__51; // @[block_division.scala 216:53]
    two_complement_buffer__52 <= two_complement__52; // @[block_division.scala 216:53]
    two_complement_buffer__53 <= two_complement__53; // @[block_division.scala 216:53]
    two_complement_buffer__54 <= two_complement__54; // @[block_division.scala 216:53]
    two_complement_buffer__55 <= two_complement__55; // @[block_division.scala 216:53]
    two_complement_buffer__56 <= two_complement__56; // @[block_division.scala 216:53]
    two_complement_buffer__57 <= two_complement__57; // @[block_division.scala 216:53]
    two_complement_buffer__58 <= two_complement__58; // @[block_division.scala 216:53]
    two_complement_buffer__59 <= two_complement__59; // @[block_division.scala 216:53]
    two_complement_buffer__60 <= two_complement__60; // @[block_division.scala 216:53]
    two_complement_buffer__61 <= two_complement__61; // @[block_division.scala 216:53]
    two_complement_buffer__62 <= two_complement__62; // @[block_division.scala 216:53]
    two_complement_buffer__63 <= two_complement__63; // @[block_division.scala 216:53]
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg <= io_man_a_0; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg <= io_sign_a_0; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_1 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_1 <= io_man_a_1; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_1 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_1 <= io_sign_a_1; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_2 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_2 <= io_man_a_2; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_2 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_2 <= io_sign_a_2; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_3 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_3 <= io_man_a_3; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_3 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_3 <= io_sign_a_3; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_4 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_4 <= io_man_a_4; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_4 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_4 <= io_sign_a_4; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_5 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_5 <= io_man_a_5; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_5 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_5 <= io_sign_a_5; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_6 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_6 <= io_man_a_6; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_6 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_6 <= io_sign_a_6; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_7 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_7 <= io_man_a_7; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_7 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_7 <= io_sign_a_7; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_8 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_8 <= io_man_a_8; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_8 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_8 <= io_sign_a_8; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_9 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_9 <= io_man_a_9; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_9 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_9 <= io_sign_a_9; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_10 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_10 <= io_man_a_10; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_10 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_10 <= io_sign_a_10; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_11 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_11 <= io_man_a_11; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_11 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_11 <= io_sign_a_11; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_12 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_12 <= io_man_a_12; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_12 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_12 <= io_sign_a_12; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_13 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_13 <= io_man_a_13; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_13 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_13 <= io_sign_a_13; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_14 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_14 <= io_man_a_14; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_14 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_14 <= io_sign_a_14; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_15 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_15 <= io_man_a_15; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_15 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_15 <= io_sign_a_15; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_16 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_16 <= io_man_a_16; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_16 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_16 <= io_sign_a_16; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_17 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_17 <= io_man_a_17; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_17 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_17 <= io_sign_a_17; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_18 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_18 <= io_man_a_18; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_18 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_18 <= io_sign_a_18; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_19 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_19 <= io_man_a_19; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_19 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_19 <= io_sign_a_19; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_20 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_20 <= io_man_a_20; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_20 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_20 <= io_sign_a_20; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_21 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_21 <= io_man_a_21; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_21 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_21 <= io_sign_a_21; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_22 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_22 <= io_man_a_22; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_22 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_22 <= io_sign_a_22; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_23 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_23 <= io_man_a_23; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_23 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_23 <= io_sign_a_23; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_24 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_24 <= io_man_a_24; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_24 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_24 <= io_sign_a_24; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_25 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_25 <= io_man_a_25; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_25 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_25 <= io_sign_a_25; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_26 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_26 <= io_man_a_26; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_26 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_26 <= io_sign_a_26; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_27 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_27 <= io_man_a_27; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_27 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_27 <= io_sign_a_27; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_28 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_28 <= io_man_a_28; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_28 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_28 <= io_sign_a_28; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_29 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_29 <= io_man_a_29; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_29 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_29 <= io_sign_a_29; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_30 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_30 <= io_man_a_30; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_30 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_30 <= io_sign_a_30; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_31 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_31 <= io_man_a_31; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_31 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_31 <= io_sign_a_31; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_32 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_32 <= io_man_a_32; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_32 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_32 <= io_sign_a_32; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_33 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_33 <= io_man_a_33; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_33 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_33 <= io_sign_a_33; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_34 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_34 <= io_man_a_34; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_34 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_34 <= io_sign_a_34; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_35 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_35 <= io_man_a_35; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_35 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_35 <= io_sign_a_35; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_36 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_36 <= io_man_a_36; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_36 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_36 <= io_sign_a_36; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_37 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_37 <= io_man_a_37; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_37 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_37 <= io_sign_a_37; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_38 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_38 <= io_man_a_38; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_38 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_38 <= io_sign_a_38; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_39 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_39 <= io_man_a_39; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_39 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_39 <= io_sign_a_39; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_40 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_40 <= io_man_a_40; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_40 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_40 <= io_sign_a_40; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_41 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_41 <= io_man_a_41; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_41 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_41 <= io_sign_a_41; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_42 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_42 <= io_man_a_42; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_42 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_42 <= io_sign_a_42; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_43 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_43 <= io_man_a_43; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_43 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_43 <= io_sign_a_43; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_44 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_44 <= io_man_a_44; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_44 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_44 <= io_sign_a_44; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_45 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_45 <= io_man_a_45; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_45 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_45 <= io_sign_a_45; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_46 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_46 <= io_man_a_46; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_46 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_46 <= io_sign_a_46; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_47 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_47 <= io_man_a_47; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_47 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_47 <= io_sign_a_47; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_48 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_48 <= io_man_a_48; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_48 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_48 <= io_sign_a_48; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_49 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_49 <= io_man_a_49; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_49 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_49 <= io_sign_a_49; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_50 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_50 <= io_man_a_50; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_50 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_50 <= io_sign_a_50; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_51 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_51 <= io_man_a_51; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_51 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_51 <= io_sign_a_51; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_52 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_52 <= io_man_a_52; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_52 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_52 <= io_sign_a_52; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_53 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_53 <= io_man_a_53; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_53 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_53 <= io_sign_a_53; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_54 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_54 <= io_man_a_54; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_54 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_54 <= io_sign_a_54; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_55 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_55 <= io_man_a_55; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_55 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_55 <= io_sign_a_55; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_56 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_56 <= io_man_a_56; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_56 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_56 <= io_sign_a_56; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_57 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_57 <= io_man_a_57; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_57 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_57 <= io_sign_a_57; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_58 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_58 <= io_man_a_58; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_58 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_58 <= io_sign_a_58; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_59 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_59 <= io_man_a_59; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_59 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_59 <= io_sign_a_59; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_60 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_60 <= io_man_a_60; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_60 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_60 <= io_sign_a_60; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_61 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_61 <= io_man_a_61; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_61 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_61 <= io_sign_a_61; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_62 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_62 <= io_man_a_62; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_62 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_62 <= io_sign_a_62; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_63 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_63 <= io_man_a_63; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_63 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_63 <= io_sign_a_63; // @[block_division.scala 206:15]
    end
    dotProductRegs_1_0 <= _dotProductRegs_0_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_1 <= _dotProductRegs_1_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_2 <= _dotProductRegs_2_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_3 <= _dotProductRegs_3_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_4 <= _dotProductRegs_4_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_5 <= _dotProductRegs_5_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_6 <= _dotProductRegs_6_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_7 <= _dotProductRegs_7_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_8 <= _dotProductRegs_8_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_9 <= _dotProductRegs_9_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_10 <= _dotProductRegs_10_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_11 <= _dotProductRegs_11_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_12 <= _dotProductRegs_12_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_13 <= _dotProductRegs_13_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_14 <= _dotProductRegs_14_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_15 <= _dotProductRegs_15_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_16 <= _dotProductRegs_16_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_17 <= _dotProductRegs_17_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_18 <= _dotProductRegs_18_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_19 <= _dotProductRegs_19_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_20 <= _dotProductRegs_20_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_21 <= _dotProductRegs_21_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_22 <= _dotProductRegs_22_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_23 <= _dotProductRegs_23_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_24 <= _dotProductRegs_24_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_25 <= _dotProductRegs_25_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_26 <= _dotProductRegs_26_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_27 <= _dotProductRegs_27_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_28 <= _dotProductRegs_28_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_29 <= _dotProductRegs_29_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_30 <= _dotProductRegs_30_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_31 <= _dotProductRegs_31_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_32 <= _dotProductRegs_32_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_33 <= _dotProductRegs_33_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_34 <= _dotProductRegs_34_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_35 <= _dotProductRegs_35_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_36 <= _dotProductRegs_36_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_37 <= _dotProductRegs_37_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_38 <= _dotProductRegs_38_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_39 <= _dotProductRegs_39_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_40 <= _dotProductRegs_40_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_41 <= _dotProductRegs_41_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_42 <= _dotProductRegs_42_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_43 <= _dotProductRegs_43_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_44 <= _dotProductRegs_44_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_45 <= _dotProductRegs_45_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_46 <= _dotProductRegs_46_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_47 <= _dotProductRegs_47_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_48 <= _dotProductRegs_48_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_49 <= _dotProductRegs_49_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_50 <= _dotProductRegs_50_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_51 <= _dotProductRegs_51_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_52 <= _dotProductRegs_52_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_53 <= _dotProductRegs_53_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_54 <= _dotProductRegs_54_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_55 <= _dotProductRegs_55_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_56 <= _dotProductRegs_56_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_57 <= _dotProductRegs_57_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_58 <= _dotProductRegs_58_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_59 <= _dotProductRegs_59_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_60 <= _dotProductRegs_60_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_61 <= _dotProductRegs_61_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_62 <= _dotProductRegs_62_T_11[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_1_63 <= _dotProductRegs_63_T_11[4:0]; // @[block_division.scala 209:25]
    signs_1_0 <= signReg_64 ^ io_sign_b_64; // @[block_division.scala 210:27]
    signs_1_1 <= signReg_65 ^ io_sign_b_65; // @[block_division.scala 210:27]
    signs_1_2 <= signReg_66 ^ io_sign_b_66; // @[block_division.scala 210:27]
    signs_1_3 <= signReg_67 ^ io_sign_b_67; // @[block_division.scala 210:27]
    signs_1_4 <= signReg_68 ^ io_sign_b_68; // @[block_division.scala 210:27]
    signs_1_5 <= signReg_69 ^ io_sign_b_69; // @[block_division.scala 210:27]
    signs_1_6 <= signReg_70 ^ io_sign_b_70; // @[block_division.scala 210:27]
    signs_1_7 <= signReg_71 ^ io_sign_b_71; // @[block_division.scala 210:27]
    signs_1_8 <= signReg_72 ^ io_sign_b_72; // @[block_division.scala 210:27]
    signs_1_9 <= signReg_73 ^ io_sign_b_73; // @[block_division.scala 210:27]
    signs_1_10 <= signReg_74 ^ io_sign_b_74; // @[block_division.scala 210:27]
    signs_1_11 <= signReg_75 ^ io_sign_b_75; // @[block_division.scala 210:27]
    signs_1_12 <= signReg_76 ^ io_sign_b_76; // @[block_division.scala 210:27]
    signs_1_13 <= signReg_77 ^ io_sign_b_77; // @[block_division.scala 210:27]
    signs_1_14 <= signReg_78 ^ io_sign_b_78; // @[block_division.scala 210:27]
    signs_1_15 <= signReg_79 ^ io_sign_b_79; // @[block_division.scala 210:27]
    signs_1_16 <= signReg_80 ^ io_sign_b_80; // @[block_division.scala 210:27]
    signs_1_17 <= signReg_81 ^ io_sign_b_81; // @[block_division.scala 210:27]
    signs_1_18 <= signReg_82 ^ io_sign_b_82; // @[block_division.scala 210:27]
    signs_1_19 <= signReg_83 ^ io_sign_b_83; // @[block_division.scala 210:27]
    signs_1_20 <= signReg_84 ^ io_sign_b_84; // @[block_division.scala 210:27]
    signs_1_21 <= signReg_85 ^ io_sign_b_85; // @[block_division.scala 210:27]
    signs_1_22 <= signReg_86 ^ io_sign_b_86; // @[block_division.scala 210:27]
    signs_1_23 <= signReg_87 ^ io_sign_b_87; // @[block_division.scala 210:27]
    signs_1_24 <= signReg_88 ^ io_sign_b_88; // @[block_division.scala 210:27]
    signs_1_25 <= signReg_89 ^ io_sign_b_89; // @[block_division.scala 210:27]
    signs_1_26 <= signReg_90 ^ io_sign_b_90; // @[block_division.scala 210:27]
    signs_1_27 <= signReg_91 ^ io_sign_b_91; // @[block_division.scala 210:27]
    signs_1_28 <= signReg_92 ^ io_sign_b_92; // @[block_division.scala 210:27]
    signs_1_29 <= signReg_93 ^ io_sign_b_93; // @[block_division.scala 210:27]
    signs_1_30 <= signReg_94 ^ io_sign_b_94; // @[block_division.scala 210:27]
    signs_1_31 <= signReg_95 ^ io_sign_b_95; // @[block_division.scala 210:27]
    signs_1_32 <= signReg_96 ^ io_sign_b_96; // @[block_division.scala 210:27]
    signs_1_33 <= signReg_97 ^ io_sign_b_97; // @[block_division.scala 210:27]
    signs_1_34 <= signReg_98 ^ io_sign_b_98; // @[block_division.scala 210:27]
    signs_1_35 <= signReg_99 ^ io_sign_b_99; // @[block_division.scala 210:27]
    signs_1_36 <= signReg_100 ^ io_sign_b_100; // @[block_division.scala 210:27]
    signs_1_37 <= signReg_101 ^ io_sign_b_101; // @[block_division.scala 210:27]
    signs_1_38 <= signReg_102 ^ io_sign_b_102; // @[block_division.scala 210:27]
    signs_1_39 <= signReg_103 ^ io_sign_b_103; // @[block_division.scala 210:27]
    signs_1_40 <= signReg_104 ^ io_sign_b_104; // @[block_division.scala 210:27]
    signs_1_41 <= signReg_105 ^ io_sign_b_105; // @[block_division.scala 210:27]
    signs_1_42 <= signReg_106 ^ io_sign_b_106; // @[block_division.scala 210:27]
    signs_1_43 <= signReg_107 ^ io_sign_b_107; // @[block_division.scala 210:27]
    signs_1_44 <= signReg_108 ^ io_sign_b_108; // @[block_division.scala 210:27]
    signs_1_45 <= signReg_109 ^ io_sign_b_109; // @[block_division.scala 210:27]
    signs_1_46 <= signReg_110 ^ io_sign_b_110; // @[block_division.scala 210:27]
    signs_1_47 <= signReg_111 ^ io_sign_b_111; // @[block_division.scala 210:27]
    signs_1_48 <= signReg_112 ^ io_sign_b_112; // @[block_division.scala 210:27]
    signs_1_49 <= signReg_113 ^ io_sign_b_113; // @[block_division.scala 210:27]
    signs_1_50 <= signReg_114 ^ io_sign_b_114; // @[block_division.scala 210:27]
    signs_1_51 <= signReg_115 ^ io_sign_b_115; // @[block_division.scala 210:27]
    signs_1_52 <= signReg_116 ^ io_sign_b_116; // @[block_division.scala 210:27]
    signs_1_53 <= signReg_117 ^ io_sign_b_117; // @[block_division.scala 210:27]
    signs_1_54 <= signReg_118 ^ io_sign_b_118; // @[block_division.scala 210:27]
    signs_1_55 <= signReg_119 ^ io_sign_b_119; // @[block_division.scala 210:27]
    signs_1_56 <= signReg_120 ^ io_sign_b_120; // @[block_division.scala 210:27]
    signs_1_57 <= signReg_121 ^ io_sign_b_121; // @[block_division.scala 210:27]
    signs_1_58 <= signReg_122 ^ io_sign_b_122; // @[block_division.scala 210:27]
    signs_1_59 <= signReg_123 ^ io_sign_b_123; // @[block_division.scala 210:27]
    signs_1_60 <= signReg_124 ^ io_sign_b_124; // @[block_division.scala 210:27]
    signs_1_61 <= signReg_125 ^ io_sign_b_125; // @[block_division.scala 210:27]
    signs_1_62 <= signReg_126 ^ io_sign_b_126; // @[block_division.scala 210:27]
    signs_1_63 <= signReg_127 ^ io_sign_b_127; // @[block_division.scala 210:27]
    if (signs_1_0) begin // @[block_division.scala 211:31]
      two_complement_1_0 <= _two_complement_0_T_11;
    end else begin
      two_complement_1_0 <= _two_complement_0_T_8;
    end
    if (signs_1_1) begin // @[block_division.scala 211:31]
      two_complement_1_1 <= _two_complement_1_T_11;
    end else begin
      two_complement_1_1 <= _two_complement_1_T_8;
    end
    if (signs_1_2) begin // @[block_division.scala 211:31]
      two_complement_1_2 <= _two_complement_2_T_11;
    end else begin
      two_complement_1_2 <= _two_complement_2_T_8;
    end
    if (signs_1_3) begin // @[block_division.scala 211:31]
      two_complement_1_3 <= _two_complement_3_T_11;
    end else begin
      two_complement_1_3 <= _two_complement_3_T_8;
    end
    if (signs_1_4) begin // @[block_division.scala 211:31]
      two_complement_1_4 <= _two_complement_4_T_11;
    end else begin
      two_complement_1_4 <= _two_complement_4_T_8;
    end
    if (signs_1_5) begin // @[block_division.scala 211:31]
      two_complement_1_5 <= _two_complement_5_T_11;
    end else begin
      two_complement_1_5 <= _two_complement_5_T_8;
    end
    if (signs_1_6) begin // @[block_division.scala 211:31]
      two_complement_1_6 <= _two_complement_6_T_11;
    end else begin
      two_complement_1_6 <= _two_complement_6_T_8;
    end
    if (signs_1_7) begin // @[block_division.scala 211:31]
      two_complement_1_7 <= _two_complement_7_T_11;
    end else begin
      two_complement_1_7 <= _two_complement_7_T_8;
    end
    if (signs_1_8) begin // @[block_division.scala 211:31]
      two_complement_1_8 <= _two_complement_8_T_11;
    end else begin
      two_complement_1_8 <= _two_complement_8_T_8;
    end
    if (signs_1_9) begin // @[block_division.scala 211:31]
      two_complement_1_9 <= _two_complement_9_T_11;
    end else begin
      two_complement_1_9 <= _two_complement_9_T_8;
    end
    if (signs_1_10) begin // @[block_division.scala 211:31]
      two_complement_1_10 <= _two_complement_10_T_11;
    end else begin
      two_complement_1_10 <= _two_complement_10_T_8;
    end
    if (signs_1_11) begin // @[block_division.scala 211:31]
      two_complement_1_11 <= _two_complement_11_T_11;
    end else begin
      two_complement_1_11 <= _two_complement_11_T_8;
    end
    if (signs_1_12) begin // @[block_division.scala 211:31]
      two_complement_1_12 <= _two_complement_12_T_11;
    end else begin
      two_complement_1_12 <= _two_complement_12_T_8;
    end
    if (signs_1_13) begin // @[block_division.scala 211:31]
      two_complement_1_13 <= _two_complement_13_T_11;
    end else begin
      two_complement_1_13 <= _two_complement_13_T_8;
    end
    if (signs_1_14) begin // @[block_division.scala 211:31]
      two_complement_1_14 <= _two_complement_14_T_11;
    end else begin
      two_complement_1_14 <= _two_complement_14_T_8;
    end
    if (signs_1_15) begin // @[block_division.scala 211:31]
      two_complement_1_15 <= _two_complement_15_T_11;
    end else begin
      two_complement_1_15 <= _two_complement_15_T_8;
    end
    if (signs_1_16) begin // @[block_division.scala 211:31]
      two_complement_1_16 <= _two_complement_16_T_11;
    end else begin
      two_complement_1_16 <= _two_complement_16_T_8;
    end
    if (signs_1_17) begin // @[block_division.scala 211:31]
      two_complement_1_17 <= _two_complement_17_T_11;
    end else begin
      two_complement_1_17 <= _two_complement_17_T_8;
    end
    if (signs_1_18) begin // @[block_division.scala 211:31]
      two_complement_1_18 <= _two_complement_18_T_11;
    end else begin
      two_complement_1_18 <= _two_complement_18_T_8;
    end
    if (signs_1_19) begin // @[block_division.scala 211:31]
      two_complement_1_19 <= _two_complement_19_T_11;
    end else begin
      two_complement_1_19 <= _two_complement_19_T_8;
    end
    if (signs_1_20) begin // @[block_division.scala 211:31]
      two_complement_1_20 <= _two_complement_20_T_11;
    end else begin
      two_complement_1_20 <= _two_complement_20_T_8;
    end
    if (signs_1_21) begin // @[block_division.scala 211:31]
      two_complement_1_21 <= _two_complement_21_T_11;
    end else begin
      two_complement_1_21 <= _two_complement_21_T_8;
    end
    if (signs_1_22) begin // @[block_division.scala 211:31]
      two_complement_1_22 <= _two_complement_22_T_11;
    end else begin
      two_complement_1_22 <= _two_complement_22_T_8;
    end
    if (signs_1_23) begin // @[block_division.scala 211:31]
      two_complement_1_23 <= _two_complement_23_T_11;
    end else begin
      two_complement_1_23 <= _two_complement_23_T_8;
    end
    if (signs_1_24) begin // @[block_division.scala 211:31]
      two_complement_1_24 <= _two_complement_24_T_11;
    end else begin
      two_complement_1_24 <= _two_complement_24_T_8;
    end
    if (signs_1_25) begin // @[block_division.scala 211:31]
      two_complement_1_25 <= _two_complement_25_T_11;
    end else begin
      two_complement_1_25 <= _two_complement_25_T_8;
    end
    if (signs_1_26) begin // @[block_division.scala 211:31]
      two_complement_1_26 <= _two_complement_26_T_11;
    end else begin
      two_complement_1_26 <= _two_complement_26_T_8;
    end
    if (signs_1_27) begin // @[block_division.scala 211:31]
      two_complement_1_27 <= _two_complement_27_T_11;
    end else begin
      two_complement_1_27 <= _two_complement_27_T_8;
    end
    if (signs_1_28) begin // @[block_division.scala 211:31]
      two_complement_1_28 <= _two_complement_28_T_11;
    end else begin
      two_complement_1_28 <= _two_complement_28_T_8;
    end
    if (signs_1_29) begin // @[block_division.scala 211:31]
      two_complement_1_29 <= _two_complement_29_T_11;
    end else begin
      two_complement_1_29 <= _two_complement_29_T_8;
    end
    if (signs_1_30) begin // @[block_division.scala 211:31]
      two_complement_1_30 <= _two_complement_30_T_11;
    end else begin
      two_complement_1_30 <= _two_complement_30_T_8;
    end
    if (signs_1_31) begin // @[block_division.scala 211:31]
      two_complement_1_31 <= _two_complement_31_T_11;
    end else begin
      two_complement_1_31 <= _two_complement_31_T_8;
    end
    if (signs_1_32) begin // @[block_division.scala 211:31]
      two_complement_1_32 <= _two_complement_32_T_11;
    end else begin
      two_complement_1_32 <= _two_complement_32_T_8;
    end
    if (signs_1_33) begin // @[block_division.scala 211:31]
      two_complement_1_33 <= _two_complement_33_T_11;
    end else begin
      two_complement_1_33 <= _two_complement_33_T_8;
    end
    if (signs_1_34) begin // @[block_division.scala 211:31]
      two_complement_1_34 <= _two_complement_34_T_11;
    end else begin
      two_complement_1_34 <= _two_complement_34_T_8;
    end
    if (signs_1_35) begin // @[block_division.scala 211:31]
      two_complement_1_35 <= _two_complement_35_T_11;
    end else begin
      two_complement_1_35 <= _two_complement_35_T_8;
    end
    if (signs_1_36) begin // @[block_division.scala 211:31]
      two_complement_1_36 <= _two_complement_36_T_11;
    end else begin
      two_complement_1_36 <= _two_complement_36_T_8;
    end
    if (signs_1_37) begin // @[block_division.scala 211:31]
      two_complement_1_37 <= _two_complement_37_T_11;
    end else begin
      two_complement_1_37 <= _two_complement_37_T_8;
    end
    if (signs_1_38) begin // @[block_division.scala 211:31]
      two_complement_1_38 <= _two_complement_38_T_11;
    end else begin
      two_complement_1_38 <= _two_complement_38_T_8;
    end
    if (signs_1_39) begin // @[block_division.scala 211:31]
      two_complement_1_39 <= _two_complement_39_T_11;
    end else begin
      two_complement_1_39 <= _two_complement_39_T_8;
    end
    if (signs_1_40) begin // @[block_division.scala 211:31]
      two_complement_1_40 <= _two_complement_40_T_11;
    end else begin
      two_complement_1_40 <= _two_complement_40_T_8;
    end
    if (signs_1_41) begin // @[block_division.scala 211:31]
      two_complement_1_41 <= _two_complement_41_T_11;
    end else begin
      two_complement_1_41 <= _two_complement_41_T_8;
    end
    if (signs_1_42) begin // @[block_division.scala 211:31]
      two_complement_1_42 <= _two_complement_42_T_11;
    end else begin
      two_complement_1_42 <= _two_complement_42_T_8;
    end
    if (signs_1_43) begin // @[block_division.scala 211:31]
      two_complement_1_43 <= _two_complement_43_T_11;
    end else begin
      two_complement_1_43 <= _two_complement_43_T_8;
    end
    if (signs_1_44) begin // @[block_division.scala 211:31]
      two_complement_1_44 <= _two_complement_44_T_11;
    end else begin
      two_complement_1_44 <= _two_complement_44_T_8;
    end
    if (signs_1_45) begin // @[block_division.scala 211:31]
      two_complement_1_45 <= _two_complement_45_T_11;
    end else begin
      two_complement_1_45 <= _two_complement_45_T_8;
    end
    if (signs_1_46) begin // @[block_division.scala 211:31]
      two_complement_1_46 <= _two_complement_46_T_11;
    end else begin
      two_complement_1_46 <= _two_complement_46_T_8;
    end
    if (signs_1_47) begin // @[block_division.scala 211:31]
      two_complement_1_47 <= _two_complement_47_T_11;
    end else begin
      two_complement_1_47 <= _two_complement_47_T_8;
    end
    if (signs_1_48) begin // @[block_division.scala 211:31]
      two_complement_1_48 <= _two_complement_48_T_11;
    end else begin
      two_complement_1_48 <= _two_complement_48_T_8;
    end
    if (signs_1_49) begin // @[block_division.scala 211:31]
      two_complement_1_49 <= _two_complement_49_T_11;
    end else begin
      two_complement_1_49 <= _two_complement_49_T_8;
    end
    if (signs_1_50) begin // @[block_division.scala 211:31]
      two_complement_1_50 <= _two_complement_50_T_11;
    end else begin
      two_complement_1_50 <= _two_complement_50_T_8;
    end
    if (signs_1_51) begin // @[block_division.scala 211:31]
      two_complement_1_51 <= _two_complement_51_T_11;
    end else begin
      two_complement_1_51 <= _two_complement_51_T_8;
    end
    if (signs_1_52) begin // @[block_division.scala 211:31]
      two_complement_1_52 <= _two_complement_52_T_11;
    end else begin
      two_complement_1_52 <= _two_complement_52_T_8;
    end
    if (signs_1_53) begin // @[block_division.scala 211:31]
      two_complement_1_53 <= _two_complement_53_T_11;
    end else begin
      two_complement_1_53 <= _two_complement_53_T_8;
    end
    if (signs_1_54) begin // @[block_division.scala 211:31]
      two_complement_1_54 <= _two_complement_54_T_11;
    end else begin
      two_complement_1_54 <= _two_complement_54_T_8;
    end
    if (signs_1_55) begin // @[block_division.scala 211:31]
      two_complement_1_55 <= _two_complement_55_T_11;
    end else begin
      two_complement_1_55 <= _two_complement_55_T_8;
    end
    if (signs_1_56) begin // @[block_division.scala 211:31]
      two_complement_1_56 <= _two_complement_56_T_11;
    end else begin
      two_complement_1_56 <= _two_complement_56_T_8;
    end
    if (signs_1_57) begin // @[block_division.scala 211:31]
      two_complement_1_57 <= _two_complement_57_T_11;
    end else begin
      two_complement_1_57 <= _two_complement_57_T_8;
    end
    if (signs_1_58) begin // @[block_division.scala 211:31]
      two_complement_1_58 <= _two_complement_58_T_11;
    end else begin
      two_complement_1_58 <= _two_complement_58_T_8;
    end
    if (signs_1_59) begin // @[block_division.scala 211:31]
      two_complement_1_59 <= _two_complement_59_T_11;
    end else begin
      two_complement_1_59 <= _two_complement_59_T_8;
    end
    if (signs_1_60) begin // @[block_division.scala 211:31]
      two_complement_1_60 <= _two_complement_60_T_11;
    end else begin
      two_complement_1_60 <= _two_complement_60_T_8;
    end
    if (signs_1_61) begin // @[block_division.scala 211:31]
      two_complement_1_61 <= _two_complement_61_T_11;
    end else begin
      two_complement_1_61 <= _two_complement_61_T_8;
    end
    if (signs_1_62) begin // @[block_division.scala 211:31]
      two_complement_1_62 <= _two_complement_62_T_11;
    end else begin
      two_complement_1_62 <= _two_complement_62_T_8;
    end
    if (signs_1_63) begin // @[block_division.scala 211:31]
      two_complement_1_63 <= _two_complement_63_T_11;
    end else begin
      two_complement_1_63 <= _two_complement_63_T_8;
    end
    two_complement_buffer_1_0 <= two_complement_1_0; // @[block_division.scala 216:53]
    two_complement_buffer_1_1 <= two_complement_1_1; // @[block_division.scala 216:53]
    two_complement_buffer_1_2 <= two_complement_1_2; // @[block_division.scala 216:53]
    two_complement_buffer_1_3 <= two_complement_1_3; // @[block_division.scala 216:53]
    two_complement_buffer_1_4 <= two_complement_1_4; // @[block_division.scala 216:53]
    two_complement_buffer_1_5 <= two_complement_1_5; // @[block_division.scala 216:53]
    two_complement_buffer_1_6 <= two_complement_1_6; // @[block_division.scala 216:53]
    two_complement_buffer_1_7 <= two_complement_1_7; // @[block_division.scala 216:53]
    two_complement_buffer_1_8 <= two_complement_1_8; // @[block_division.scala 216:53]
    two_complement_buffer_1_9 <= two_complement_1_9; // @[block_division.scala 216:53]
    two_complement_buffer_1_10 <= two_complement_1_10; // @[block_division.scala 216:53]
    two_complement_buffer_1_11 <= two_complement_1_11; // @[block_division.scala 216:53]
    two_complement_buffer_1_12 <= two_complement_1_12; // @[block_division.scala 216:53]
    two_complement_buffer_1_13 <= two_complement_1_13; // @[block_division.scala 216:53]
    two_complement_buffer_1_14 <= two_complement_1_14; // @[block_division.scala 216:53]
    two_complement_buffer_1_15 <= two_complement_1_15; // @[block_division.scala 216:53]
    two_complement_buffer_1_16 <= two_complement_1_16; // @[block_division.scala 216:53]
    two_complement_buffer_1_17 <= two_complement_1_17; // @[block_division.scala 216:53]
    two_complement_buffer_1_18 <= two_complement_1_18; // @[block_division.scala 216:53]
    two_complement_buffer_1_19 <= two_complement_1_19; // @[block_division.scala 216:53]
    two_complement_buffer_1_20 <= two_complement_1_20; // @[block_division.scala 216:53]
    two_complement_buffer_1_21 <= two_complement_1_21; // @[block_division.scala 216:53]
    two_complement_buffer_1_22 <= two_complement_1_22; // @[block_division.scala 216:53]
    two_complement_buffer_1_23 <= two_complement_1_23; // @[block_division.scala 216:53]
    two_complement_buffer_1_24 <= two_complement_1_24; // @[block_division.scala 216:53]
    two_complement_buffer_1_25 <= two_complement_1_25; // @[block_division.scala 216:53]
    two_complement_buffer_1_26 <= two_complement_1_26; // @[block_division.scala 216:53]
    two_complement_buffer_1_27 <= two_complement_1_27; // @[block_division.scala 216:53]
    two_complement_buffer_1_28 <= two_complement_1_28; // @[block_division.scala 216:53]
    two_complement_buffer_1_29 <= two_complement_1_29; // @[block_division.scala 216:53]
    two_complement_buffer_1_30 <= two_complement_1_30; // @[block_division.scala 216:53]
    two_complement_buffer_1_31 <= two_complement_1_31; // @[block_division.scala 216:53]
    two_complement_buffer_1_32 <= two_complement_1_32; // @[block_division.scala 216:53]
    two_complement_buffer_1_33 <= two_complement_1_33; // @[block_division.scala 216:53]
    two_complement_buffer_1_34 <= two_complement_1_34; // @[block_division.scala 216:53]
    two_complement_buffer_1_35 <= two_complement_1_35; // @[block_division.scala 216:53]
    two_complement_buffer_1_36 <= two_complement_1_36; // @[block_division.scala 216:53]
    two_complement_buffer_1_37 <= two_complement_1_37; // @[block_division.scala 216:53]
    two_complement_buffer_1_38 <= two_complement_1_38; // @[block_division.scala 216:53]
    two_complement_buffer_1_39 <= two_complement_1_39; // @[block_division.scala 216:53]
    two_complement_buffer_1_40 <= two_complement_1_40; // @[block_division.scala 216:53]
    two_complement_buffer_1_41 <= two_complement_1_41; // @[block_division.scala 216:53]
    two_complement_buffer_1_42 <= two_complement_1_42; // @[block_division.scala 216:53]
    two_complement_buffer_1_43 <= two_complement_1_43; // @[block_division.scala 216:53]
    two_complement_buffer_1_44 <= two_complement_1_44; // @[block_division.scala 216:53]
    two_complement_buffer_1_45 <= two_complement_1_45; // @[block_division.scala 216:53]
    two_complement_buffer_1_46 <= two_complement_1_46; // @[block_division.scala 216:53]
    two_complement_buffer_1_47 <= two_complement_1_47; // @[block_division.scala 216:53]
    two_complement_buffer_1_48 <= two_complement_1_48; // @[block_division.scala 216:53]
    two_complement_buffer_1_49 <= two_complement_1_49; // @[block_division.scala 216:53]
    two_complement_buffer_1_50 <= two_complement_1_50; // @[block_division.scala 216:53]
    two_complement_buffer_1_51 <= two_complement_1_51; // @[block_division.scala 216:53]
    two_complement_buffer_1_52 <= two_complement_1_52; // @[block_division.scala 216:53]
    two_complement_buffer_1_53 <= two_complement_1_53; // @[block_division.scala 216:53]
    two_complement_buffer_1_54 <= two_complement_1_54; // @[block_division.scala 216:53]
    two_complement_buffer_1_55 <= two_complement_1_55; // @[block_division.scala 216:53]
    two_complement_buffer_1_56 <= two_complement_1_56; // @[block_division.scala 216:53]
    two_complement_buffer_1_57 <= two_complement_1_57; // @[block_division.scala 216:53]
    two_complement_buffer_1_58 <= two_complement_1_58; // @[block_division.scala 216:53]
    two_complement_buffer_1_59 <= two_complement_1_59; // @[block_division.scala 216:53]
    two_complement_buffer_1_60 <= two_complement_1_60; // @[block_division.scala 216:53]
    two_complement_buffer_1_61 <= two_complement_1_61; // @[block_division.scala 216:53]
    two_complement_buffer_1_62 <= two_complement_1_62; // @[block_division.scala 216:53]
    two_complement_buffer_1_63 <= two_complement_1_63; // @[block_division.scala 216:53]
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_64 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_64 <= io_man_a_64; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_64 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_64 <= io_sign_a_64; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_65 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_65 <= io_man_a_65; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_65 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_65 <= io_sign_a_65; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_66 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_66 <= io_man_a_66; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_66 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_66 <= io_sign_a_66; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_67 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_67 <= io_man_a_67; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_67 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_67 <= io_sign_a_67; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_68 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_68 <= io_man_a_68; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_68 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_68 <= io_sign_a_68; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_69 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_69 <= io_man_a_69; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_69 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_69 <= io_sign_a_69; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_70 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_70 <= io_man_a_70; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_70 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_70 <= io_sign_a_70; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_71 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_71 <= io_man_a_71; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_71 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_71 <= io_sign_a_71; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_72 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_72 <= io_man_a_72; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_72 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_72 <= io_sign_a_72; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_73 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_73 <= io_man_a_73; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_73 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_73 <= io_sign_a_73; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_74 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_74 <= io_man_a_74; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_74 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_74 <= io_sign_a_74; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_75 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_75 <= io_man_a_75; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_75 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_75 <= io_sign_a_75; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_76 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_76 <= io_man_a_76; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_76 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_76 <= io_sign_a_76; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_77 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_77 <= io_man_a_77; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_77 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_77 <= io_sign_a_77; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_78 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_78 <= io_man_a_78; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_78 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_78 <= io_sign_a_78; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_79 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_79 <= io_man_a_79; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_79 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_79 <= io_sign_a_79; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_80 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_80 <= io_man_a_80; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_80 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_80 <= io_sign_a_80; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_81 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_81 <= io_man_a_81; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_81 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_81 <= io_sign_a_81; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_82 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_82 <= io_man_a_82; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_82 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_82 <= io_sign_a_82; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_83 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_83 <= io_man_a_83; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_83 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_83 <= io_sign_a_83; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_84 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_84 <= io_man_a_84; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_84 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_84 <= io_sign_a_84; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_85 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_85 <= io_man_a_85; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_85 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_85 <= io_sign_a_85; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_86 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_86 <= io_man_a_86; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_86 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_86 <= io_sign_a_86; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_87 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_87 <= io_man_a_87; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_87 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_87 <= io_sign_a_87; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_88 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_88 <= io_man_a_88; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_88 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_88 <= io_sign_a_88; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_89 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_89 <= io_man_a_89; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_89 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_89 <= io_sign_a_89; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_90 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_90 <= io_man_a_90; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_90 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_90 <= io_sign_a_90; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_91 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_91 <= io_man_a_91; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_91 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_91 <= io_sign_a_91; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_92 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_92 <= io_man_a_92; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_92 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_92 <= io_sign_a_92; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_93 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_93 <= io_man_a_93; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_93 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_93 <= io_sign_a_93; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_94 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_94 <= io_man_a_94; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_94 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_94 <= io_sign_a_94; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_95 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_95 <= io_man_a_95; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_95 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_95 <= io_sign_a_95; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_96 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_96 <= io_man_a_96; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_96 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_96 <= io_sign_a_96; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_97 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_97 <= io_man_a_97; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_97 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_97 <= io_sign_a_97; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_98 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_98 <= io_man_a_98; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_98 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_98 <= io_sign_a_98; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_99 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_99 <= io_man_a_99; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_99 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_99 <= io_sign_a_99; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_100 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_100 <= io_man_a_100; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_100 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_100 <= io_sign_a_100; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_101 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_101 <= io_man_a_101; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_101 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_101 <= io_sign_a_101; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_102 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_102 <= io_man_a_102; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_102 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_102 <= io_sign_a_102; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_103 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_103 <= io_man_a_103; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_103 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_103 <= io_sign_a_103; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_104 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_104 <= io_man_a_104; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_104 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_104 <= io_sign_a_104; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_105 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_105 <= io_man_a_105; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_105 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_105 <= io_sign_a_105; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_106 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_106 <= io_man_a_106; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_106 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_106 <= io_sign_a_106; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_107 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_107 <= io_man_a_107; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_107 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_107 <= io_sign_a_107; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_108 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_108 <= io_man_a_108; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_108 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_108 <= io_sign_a_108; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_109 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_109 <= io_man_a_109; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_109 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_109 <= io_sign_a_109; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_110 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_110 <= io_man_a_110; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_110 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_110 <= io_sign_a_110; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_111 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_111 <= io_man_a_111; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_111 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_111 <= io_sign_a_111; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_112 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_112 <= io_man_a_112; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_112 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_112 <= io_sign_a_112; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_113 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_113 <= io_man_a_113; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_113 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_113 <= io_sign_a_113; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_114 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_114 <= io_man_a_114; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_114 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_114 <= io_sign_a_114; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_115 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_115 <= io_man_a_115; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_115 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_115 <= io_sign_a_115; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_116 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_116 <= io_man_a_116; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_116 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_116 <= io_sign_a_116; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_117 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_117 <= io_man_a_117; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_117 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_117 <= io_sign_a_117; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_118 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_118 <= io_man_a_118; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_118 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_118 <= io_sign_a_118; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_119 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_119 <= io_man_a_119; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_119 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_119 <= io_sign_a_119; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_120 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_120 <= io_man_a_120; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_120 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_120 <= io_sign_a_120; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_121 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_121 <= io_man_a_121; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_121 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_121 <= io_sign_a_121; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_122 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_122 <= io_man_a_122; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_122 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_122 <= io_sign_a_122; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_123 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_123 <= io_man_a_123; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_123 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_123 <= io_sign_a_123; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_124 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_124 <= io_man_a_124; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_124 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_124 <= io_sign_a_124; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_125 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_125 <= io_man_a_125; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_125 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_125 <= io_sign_a_125; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_126 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_126 <= io_man_a_126; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_126 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_126 <= io_sign_a_126; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_127 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_127 <= io_man_a_127; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_127 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_127 <= io_sign_a_127; // @[block_division.scala 206:15]
    end
    dotProductRegs_2_0 <= _dotProductRegs_0_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_1 <= _dotProductRegs_1_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_2 <= _dotProductRegs_2_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_3 <= _dotProductRegs_3_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_4 <= _dotProductRegs_4_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_5 <= _dotProductRegs_5_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_6 <= _dotProductRegs_6_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_7 <= _dotProductRegs_7_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_8 <= _dotProductRegs_8_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_9 <= _dotProductRegs_9_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_10 <= _dotProductRegs_10_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_11 <= _dotProductRegs_11_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_12 <= _dotProductRegs_12_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_13 <= _dotProductRegs_13_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_14 <= _dotProductRegs_14_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_15 <= _dotProductRegs_15_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_16 <= _dotProductRegs_16_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_17 <= _dotProductRegs_17_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_18 <= _dotProductRegs_18_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_19 <= _dotProductRegs_19_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_20 <= _dotProductRegs_20_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_21 <= _dotProductRegs_21_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_22 <= _dotProductRegs_22_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_23 <= _dotProductRegs_23_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_24 <= _dotProductRegs_24_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_25 <= _dotProductRegs_25_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_26 <= _dotProductRegs_26_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_27 <= _dotProductRegs_27_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_28 <= _dotProductRegs_28_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_29 <= _dotProductRegs_29_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_30 <= _dotProductRegs_30_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_31 <= _dotProductRegs_31_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_32 <= _dotProductRegs_32_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_33 <= _dotProductRegs_33_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_34 <= _dotProductRegs_34_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_35 <= _dotProductRegs_35_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_36 <= _dotProductRegs_36_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_37 <= _dotProductRegs_37_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_38 <= _dotProductRegs_38_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_39 <= _dotProductRegs_39_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_40 <= _dotProductRegs_40_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_41 <= _dotProductRegs_41_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_42 <= _dotProductRegs_42_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_43 <= _dotProductRegs_43_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_44 <= _dotProductRegs_44_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_45 <= _dotProductRegs_45_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_46 <= _dotProductRegs_46_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_47 <= _dotProductRegs_47_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_48 <= _dotProductRegs_48_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_49 <= _dotProductRegs_49_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_50 <= _dotProductRegs_50_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_51 <= _dotProductRegs_51_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_52 <= _dotProductRegs_52_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_53 <= _dotProductRegs_53_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_54 <= _dotProductRegs_54_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_55 <= _dotProductRegs_55_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_56 <= _dotProductRegs_56_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_57 <= _dotProductRegs_57_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_58 <= _dotProductRegs_58_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_59 <= _dotProductRegs_59_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_60 <= _dotProductRegs_60_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_61 <= _dotProductRegs_61_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_62 <= _dotProductRegs_62_T_17[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_2_63 <= _dotProductRegs_63_T_17[4:0]; // @[block_division.scala 209:25]
    signs_2_0 <= signReg_128 ^ io_sign_b_128; // @[block_division.scala 210:27]
    signs_2_1 <= signReg_129 ^ io_sign_b_129; // @[block_division.scala 210:27]
    signs_2_2 <= signReg_130 ^ io_sign_b_130; // @[block_division.scala 210:27]
    signs_2_3 <= signReg_131 ^ io_sign_b_131; // @[block_division.scala 210:27]
    signs_2_4 <= signReg_132 ^ io_sign_b_132; // @[block_division.scala 210:27]
    signs_2_5 <= signReg_133 ^ io_sign_b_133; // @[block_division.scala 210:27]
    signs_2_6 <= signReg_134 ^ io_sign_b_134; // @[block_division.scala 210:27]
    signs_2_7 <= signReg_135 ^ io_sign_b_135; // @[block_division.scala 210:27]
    signs_2_8 <= signReg_136 ^ io_sign_b_136; // @[block_division.scala 210:27]
    signs_2_9 <= signReg_137 ^ io_sign_b_137; // @[block_division.scala 210:27]
    signs_2_10 <= signReg_138 ^ io_sign_b_138; // @[block_division.scala 210:27]
    signs_2_11 <= signReg_139 ^ io_sign_b_139; // @[block_division.scala 210:27]
    signs_2_12 <= signReg_140 ^ io_sign_b_140; // @[block_division.scala 210:27]
    signs_2_13 <= signReg_141 ^ io_sign_b_141; // @[block_division.scala 210:27]
    signs_2_14 <= signReg_142 ^ io_sign_b_142; // @[block_division.scala 210:27]
    signs_2_15 <= signReg_143 ^ io_sign_b_143; // @[block_division.scala 210:27]
    signs_2_16 <= signReg_144 ^ io_sign_b_144; // @[block_division.scala 210:27]
    signs_2_17 <= signReg_145 ^ io_sign_b_145; // @[block_division.scala 210:27]
    signs_2_18 <= signReg_146 ^ io_sign_b_146; // @[block_division.scala 210:27]
    signs_2_19 <= signReg_147 ^ io_sign_b_147; // @[block_division.scala 210:27]
    signs_2_20 <= signReg_148 ^ io_sign_b_148; // @[block_division.scala 210:27]
    signs_2_21 <= signReg_149 ^ io_sign_b_149; // @[block_division.scala 210:27]
    signs_2_22 <= signReg_150 ^ io_sign_b_150; // @[block_division.scala 210:27]
    signs_2_23 <= signReg_151 ^ io_sign_b_151; // @[block_division.scala 210:27]
    signs_2_24 <= signReg_152 ^ io_sign_b_152; // @[block_division.scala 210:27]
    signs_2_25 <= signReg_153 ^ io_sign_b_153; // @[block_division.scala 210:27]
    signs_2_26 <= signReg_154 ^ io_sign_b_154; // @[block_division.scala 210:27]
    signs_2_27 <= signReg_155 ^ io_sign_b_155; // @[block_division.scala 210:27]
    signs_2_28 <= signReg_156 ^ io_sign_b_156; // @[block_division.scala 210:27]
    signs_2_29 <= signReg_157 ^ io_sign_b_157; // @[block_division.scala 210:27]
    signs_2_30 <= signReg_158 ^ io_sign_b_158; // @[block_division.scala 210:27]
    signs_2_31 <= signReg_159 ^ io_sign_b_159; // @[block_division.scala 210:27]
    signs_2_32 <= signReg_160 ^ io_sign_b_160; // @[block_division.scala 210:27]
    signs_2_33 <= signReg_161 ^ io_sign_b_161; // @[block_division.scala 210:27]
    signs_2_34 <= signReg_162 ^ io_sign_b_162; // @[block_division.scala 210:27]
    signs_2_35 <= signReg_163 ^ io_sign_b_163; // @[block_division.scala 210:27]
    signs_2_36 <= signReg_164 ^ io_sign_b_164; // @[block_division.scala 210:27]
    signs_2_37 <= signReg_165 ^ io_sign_b_165; // @[block_division.scala 210:27]
    signs_2_38 <= signReg_166 ^ io_sign_b_166; // @[block_division.scala 210:27]
    signs_2_39 <= signReg_167 ^ io_sign_b_167; // @[block_division.scala 210:27]
    signs_2_40 <= signReg_168 ^ io_sign_b_168; // @[block_division.scala 210:27]
    signs_2_41 <= signReg_169 ^ io_sign_b_169; // @[block_division.scala 210:27]
    signs_2_42 <= signReg_170 ^ io_sign_b_170; // @[block_division.scala 210:27]
    signs_2_43 <= signReg_171 ^ io_sign_b_171; // @[block_division.scala 210:27]
    signs_2_44 <= signReg_172 ^ io_sign_b_172; // @[block_division.scala 210:27]
    signs_2_45 <= signReg_173 ^ io_sign_b_173; // @[block_division.scala 210:27]
    signs_2_46 <= signReg_174 ^ io_sign_b_174; // @[block_division.scala 210:27]
    signs_2_47 <= signReg_175 ^ io_sign_b_175; // @[block_division.scala 210:27]
    signs_2_48 <= signReg_176 ^ io_sign_b_176; // @[block_division.scala 210:27]
    signs_2_49 <= signReg_177 ^ io_sign_b_177; // @[block_division.scala 210:27]
    signs_2_50 <= signReg_178 ^ io_sign_b_178; // @[block_division.scala 210:27]
    signs_2_51 <= signReg_179 ^ io_sign_b_179; // @[block_division.scala 210:27]
    signs_2_52 <= signReg_180 ^ io_sign_b_180; // @[block_division.scala 210:27]
    signs_2_53 <= signReg_181 ^ io_sign_b_181; // @[block_division.scala 210:27]
    signs_2_54 <= signReg_182 ^ io_sign_b_182; // @[block_division.scala 210:27]
    signs_2_55 <= signReg_183 ^ io_sign_b_183; // @[block_division.scala 210:27]
    signs_2_56 <= signReg_184 ^ io_sign_b_184; // @[block_division.scala 210:27]
    signs_2_57 <= signReg_185 ^ io_sign_b_185; // @[block_division.scala 210:27]
    signs_2_58 <= signReg_186 ^ io_sign_b_186; // @[block_division.scala 210:27]
    signs_2_59 <= signReg_187 ^ io_sign_b_187; // @[block_division.scala 210:27]
    signs_2_60 <= signReg_188 ^ io_sign_b_188; // @[block_division.scala 210:27]
    signs_2_61 <= signReg_189 ^ io_sign_b_189; // @[block_division.scala 210:27]
    signs_2_62 <= signReg_190 ^ io_sign_b_190; // @[block_division.scala 210:27]
    signs_2_63 <= signReg_191 ^ io_sign_b_191; // @[block_division.scala 210:27]
    if (signs_2_0) begin // @[block_division.scala 211:31]
      two_complement_2_0 <= _two_complement_0_T_18;
    end else begin
      two_complement_2_0 <= _two_complement_0_T_15;
    end
    if (signs_2_1) begin // @[block_division.scala 211:31]
      two_complement_2_1 <= _two_complement_1_T_18;
    end else begin
      two_complement_2_1 <= _two_complement_1_T_15;
    end
    if (signs_2_2) begin // @[block_division.scala 211:31]
      two_complement_2_2 <= _two_complement_2_T_18;
    end else begin
      two_complement_2_2 <= _two_complement_2_T_15;
    end
    if (signs_2_3) begin // @[block_division.scala 211:31]
      two_complement_2_3 <= _two_complement_3_T_18;
    end else begin
      two_complement_2_3 <= _two_complement_3_T_15;
    end
    if (signs_2_4) begin // @[block_division.scala 211:31]
      two_complement_2_4 <= _two_complement_4_T_18;
    end else begin
      two_complement_2_4 <= _two_complement_4_T_15;
    end
    if (signs_2_5) begin // @[block_division.scala 211:31]
      two_complement_2_5 <= _two_complement_5_T_18;
    end else begin
      two_complement_2_5 <= _two_complement_5_T_15;
    end
    if (signs_2_6) begin // @[block_division.scala 211:31]
      two_complement_2_6 <= _two_complement_6_T_18;
    end else begin
      two_complement_2_6 <= _two_complement_6_T_15;
    end
    if (signs_2_7) begin // @[block_division.scala 211:31]
      two_complement_2_7 <= _two_complement_7_T_18;
    end else begin
      two_complement_2_7 <= _two_complement_7_T_15;
    end
    if (signs_2_8) begin // @[block_division.scala 211:31]
      two_complement_2_8 <= _two_complement_8_T_18;
    end else begin
      two_complement_2_8 <= _two_complement_8_T_15;
    end
    if (signs_2_9) begin // @[block_division.scala 211:31]
      two_complement_2_9 <= _two_complement_9_T_18;
    end else begin
      two_complement_2_9 <= _two_complement_9_T_15;
    end
    if (signs_2_10) begin // @[block_division.scala 211:31]
      two_complement_2_10 <= _two_complement_10_T_18;
    end else begin
      two_complement_2_10 <= _two_complement_10_T_15;
    end
    if (signs_2_11) begin // @[block_division.scala 211:31]
      two_complement_2_11 <= _two_complement_11_T_18;
    end else begin
      two_complement_2_11 <= _two_complement_11_T_15;
    end
    if (signs_2_12) begin // @[block_division.scala 211:31]
      two_complement_2_12 <= _two_complement_12_T_18;
    end else begin
      two_complement_2_12 <= _two_complement_12_T_15;
    end
    if (signs_2_13) begin // @[block_division.scala 211:31]
      two_complement_2_13 <= _two_complement_13_T_18;
    end else begin
      two_complement_2_13 <= _two_complement_13_T_15;
    end
    if (signs_2_14) begin // @[block_division.scala 211:31]
      two_complement_2_14 <= _two_complement_14_T_18;
    end else begin
      two_complement_2_14 <= _two_complement_14_T_15;
    end
    if (signs_2_15) begin // @[block_division.scala 211:31]
      two_complement_2_15 <= _two_complement_15_T_18;
    end else begin
      two_complement_2_15 <= _two_complement_15_T_15;
    end
    if (signs_2_16) begin // @[block_division.scala 211:31]
      two_complement_2_16 <= _two_complement_16_T_18;
    end else begin
      two_complement_2_16 <= _two_complement_16_T_15;
    end
    if (signs_2_17) begin // @[block_division.scala 211:31]
      two_complement_2_17 <= _two_complement_17_T_18;
    end else begin
      two_complement_2_17 <= _two_complement_17_T_15;
    end
    if (signs_2_18) begin // @[block_division.scala 211:31]
      two_complement_2_18 <= _two_complement_18_T_18;
    end else begin
      two_complement_2_18 <= _two_complement_18_T_15;
    end
    if (signs_2_19) begin // @[block_division.scala 211:31]
      two_complement_2_19 <= _two_complement_19_T_18;
    end else begin
      two_complement_2_19 <= _two_complement_19_T_15;
    end
    if (signs_2_20) begin // @[block_division.scala 211:31]
      two_complement_2_20 <= _two_complement_20_T_18;
    end else begin
      two_complement_2_20 <= _two_complement_20_T_15;
    end
    if (signs_2_21) begin // @[block_division.scala 211:31]
      two_complement_2_21 <= _two_complement_21_T_18;
    end else begin
      two_complement_2_21 <= _two_complement_21_T_15;
    end
    if (signs_2_22) begin // @[block_division.scala 211:31]
      two_complement_2_22 <= _two_complement_22_T_18;
    end else begin
      two_complement_2_22 <= _two_complement_22_T_15;
    end
    if (signs_2_23) begin // @[block_division.scala 211:31]
      two_complement_2_23 <= _two_complement_23_T_18;
    end else begin
      two_complement_2_23 <= _two_complement_23_T_15;
    end
    if (signs_2_24) begin // @[block_division.scala 211:31]
      two_complement_2_24 <= _two_complement_24_T_18;
    end else begin
      two_complement_2_24 <= _two_complement_24_T_15;
    end
    if (signs_2_25) begin // @[block_division.scala 211:31]
      two_complement_2_25 <= _two_complement_25_T_18;
    end else begin
      two_complement_2_25 <= _two_complement_25_T_15;
    end
    if (signs_2_26) begin // @[block_division.scala 211:31]
      two_complement_2_26 <= _two_complement_26_T_18;
    end else begin
      two_complement_2_26 <= _two_complement_26_T_15;
    end
    if (signs_2_27) begin // @[block_division.scala 211:31]
      two_complement_2_27 <= _two_complement_27_T_18;
    end else begin
      two_complement_2_27 <= _two_complement_27_T_15;
    end
    if (signs_2_28) begin // @[block_division.scala 211:31]
      two_complement_2_28 <= _two_complement_28_T_18;
    end else begin
      two_complement_2_28 <= _two_complement_28_T_15;
    end
    if (signs_2_29) begin // @[block_division.scala 211:31]
      two_complement_2_29 <= _two_complement_29_T_18;
    end else begin
      two_complement_2_29 <= _two_complement_29_T_15;
    end
    if (signs_2_30) begin // @[block_division.scala 211:31]
      two_complement_2_30 <= _two_complement_30_T_18;
    end else begin
      two_complement_2_30 <= _two_complement_30_T_15;
    end
    if (signs_2_31) begin // @[block_division.scala 211:31]
      two_complement_2_31 <= _two_complement_31_T_18;
    end else begin
      two_complement_2_31 <= _two_complement_31_T_15;
    end
    if (signs_2_32) begin // @[block_division.scala 211:31]
      two_complement_2_32 <= _two_complement_32_T_18;
    end else begin
      two_complement_2_32 <= _two_complement_32_T_15;
    end
    if (signs_2_33) begin // @[block_division.scala 211:31]
      two_complement_2_33 <= _two_complement_33_T_18;
    end else begin
      two_complement_2_33 <= _two_complement_33_T_15;
    end
    if (signs_2_34) begin // @[block_division.scala 211:31]
      two_complement_2_34 <= _two_complement_34_T_18;
    end else begin
      two_complement_2_34 <= _two_complement_34_T_15;
    end
    if (signs_2_35) begin // @[block_division.scala 211:31]
      two_complement_2_35 <= _two_complement_35_T_18;
    end else begin
      two_complement_2_35 <= _two_complement_35_T_15;
    end
    if (signs_2_36) begin // @[block_division.scala 211:31]
      two_complement_2_36 <= _two_complement_36_T_18;
    end else begin
      two_complement_2_36 <= _two_complement_36_T_15;
    end
    if (signs_2_37) begin // @[block_division.scala 211:31]
      two_complement_2_37 <= _two_complement_37_T_18;
    end else begin
      two_complement_2_37 <= _two_complement_37_T_15;
    end
    if (signs_2_38) begin // @[block_division.scala 211:31]
      two_complement_2_38 <= _two_complement_38_T_18;
    end else begin
      two_complement_2_38 <= _two_complement_38_T_15;
    end
    if (signs_2_39) begin // @[block_division.scala 211:31]
      two_complement_2_39 <= _two_complement_39_T_18;
    end else begin
      two_complement_2_39 <= _two_complement_39_T_15;
    end
    if (signs_2_40) begin // @[block_division.scala 211:31]
      two_complement_2_40 <= _two_complement_40_T_18;
    end else begin
      two_complement_2_40 <= _two_complement_40_T_15;
    end
    if (signs_2_41) begin // @[block_division.scala 211:31]
      two_complement_2_41 <= _two_complement_41_T_18;
    end else begin
      two_complement_2_41 <= _two_complement_41_T_15;
    end
    if (signs_2_42) begin // @[block_division.scala 211:31]
      two_complement_2_42 <= _two_complement_42_T_18;
    end else begin
      two_complement_2_42 <= _two_complement_42_T_15;
    end
    if (signs_2_43) begin // @[block_division.scala 211:31]
      two_complement_2_43 <= _two_complement_43_T_18;
    end else begin
      two_complement_2_43 <= _two_complement_43_T_15;
    end
    if (signs_2_44) begin // @[block_division.scala 211:31]
      two_complement_2_44 <= _two_complement_44_T_18;
    end else begin
      two_complement_2_44 <= _two_complement_44_T_15;
    end
    if (signs_2_45) begin // @[block_division.scala 211:31]
      two_complement_2_45 <= _two_complement_45_T_18;
    end else begin
      two_complement_2_45 <= _two_complement_45_T_15;
    end
    if (signs_2_46) begin // @[block_division.scala 211:31]
      two_complement_2_46 <= _two_complement_46_T_18;
    end else begin
      two_complement_2_46 <= _two_complement_46_T_15;
    end
    if (signs_2_47) begin // @[block_division.scala 211:31]
      two_complement_2_47 <= _two_complement_47_T_18;
    end else begin
      two_complement_2_47 <= _two_complement_47_T_15;
    end
    if (signs_2_48) begin // @[block_division.scala 211:31]
      two_complement_2_48 <= _two_complement_48_T_18;
    end else begin
      two_complement_2_48 <= _two_complement_48_T_15;
    end
    if (signs_2_49) begin // @[block_division.scala 211:31]
      two_complement_2_49 <= _two_complement_49_T_18;
    end else begin
      two_complement_2_49 <= _two_complement_49_T_15;
    end
    if (signs_2_50) begin // @[block_division.scala 211:31]
      two_complement_2_50 <= _two_complement_50_T_18;
    end else begin
      two_complement_2_50 <= _two_complement_50_T_15;
    end
    if (signs_2_51) begin // @[block_division.scala 211:31]
      two_complement_2_51 <= _two_complement_51_T_18;
    end else begin
      two_complement_2_51 <= _two_complement_51_T_15;
    end
    if (signs_2_52) begin // @[block_division.scala 211:31]
      two_complement_2_52 <= _two_complement_52_T_18;
    end else begin
      two_complement_2_52 <= _two_complement_52_T_15;
    end
    if (signs_2_53) begin // @[block_division.scala 211:31]
      two_complement_2_53 <= _two_complement_53_T_18;
    end else begin
      two_complement_2_53 <= _two_complement_53_T_15;
    end
    if (signs_2_54) begin // @[block_division.scala 211:31]
      two_complement_2_54 <= _two_complement_54_T_18;
    end else begin
      two_complement_2_54 <= _two_complement_54_T_15;
    end
    if (signs_2_55) begin // @[block_division.scala 211:31]
      two_complement_2_55 <= _two_complement_55_T_18;
    end else begin
      two_complement_2_55 <= _two_complement_55_T_15;
    end
    if (signs_2_56) begin // @[block_division.scala 211:31]
      two_complement_2_56 <= _two_complement_56_T_18;
    end else begin
      two_complement_2_56 <= _two_complement_56_T_15;
    end
    if (signs_2_57) begin // @[block_division.scala 211:31]
      two_complement_2_57 <= _two_complement_57_T_18;
    end else begin
      two_complement_2_57 <= _two_complement_57_T_15;
    end
    if (signs_2_58) begin // @[block_division.scala 211:31]
      two_complement_2_58 <= _two_complement_58_T_18;
    end else begin
      two_complement_2_58 <= _two_complement_58_T_15;
    end
    if (signs_2_59) begin // @[block_division.scala 211:31]
      two_complement_2_59 <= _two_complement_59_T_18;
    end else begin
      two_complement_2_59 <= _two_complement_59_T_15;
    end
    if (signs_2_60) begin // @[block_division.scala 211:31]
      two_complement_2_60 <= _two_complement_60_T_18;
    end else begin
      two_complement_2_60 <= _two_complement_60_T_15;
    end
    if (signs_2_61) begin // @[block_division.scala 211:31]
      two_complement_2_61 <= _two_complement_61_T_18;
    end else begin
      two_complement_2_61 <= _two_complement_61_T_15;
    end
    if (signs_2_62) begin // @[block_division.scala 211:31]
      two_complement_2_62 <= _two_complement_62_T_18;
    end else begin
      two_complement_2_62 <= _two_complement_62_T_15;
    end
    if (signs_2_63) begin // @[block_division.scala 211:31]
      two_complement_2_63 <= _two_complement_63_T_18;
    end else begin
      two_complement_2_63 <= _two_complement_63_T_15;
    end
    two_complement_buffer_2_0 <= two_complement_2_0; // @[block_division.scala 216:53]
    two_complement_buffer_2_1 <= two_complement_2_1; // @[block_division.scala 216:53]
    two_complement_buffer_2_2 <= two_complement_2_2; // @[block_division.scala 216:53]
    two_complement_buffer_2_3 <= two_complement_2_3; // @[block_division.scala 216:53]
    two_complement_buffer_2_4 <= two_complement_2_4; // @[block_division.scala 216:53]
    two_complement_buffer_2_5 <= two_complement_2_5; // @[block_division.scala 216:53]
    two_complement_buffer_2_6 <= two_complement_2_6; // @[block_division.scala 216:53]
    two_complement_buffer_2_7 <= two_complement_2_7; // @[block_division.scala 216:53]
    two_complement_buffer_2_8 <= two_complement_2_8; // @[block_division.scala 216:53]
    two_complement_buffer_2_9 <= two_complement_2_9; // @[block_division.scala 216:53]
    two_complement_buffer_2_10 <= two_complement_2_10; // @[block_division.scala 216:53]
    two_complement_buffer_2_11 <= two_complement_2_11; // @[block_division.scala 216:53]
    two_complement_buffer_2_12 <= two_complement_2_12; // @[block_division.scala 216:53]
    two_complement_buffer_2_13 <= two_complement_2_13; // @[block_division.scala 216:53]
    two_complement_buffer_2_14 <= two_complement_2_14; // @[block_division.scala 216:53]
    two_complement_buffer_2_15 <= two_complement_2_15; // @[block_division.scala 216:53]
    two_complement_buffer_2_16 <= two_complement_2_16; // @[block_division.scala 216:53]
    two_complement_buffer_2_17 <= two_complement_2_17; // @[block_division.scala 216:53]
    two_complement_buffer_2_18 <= two_complement_2_18; // @[block_division.scala 216:53]
    two_complement_buffer_2_19 <= two_complement_2_19; // @[block_division.scala 216:53]
    two_complement_buffer_2_20 <= two_complement_2_20; // @[block_division.scala 216:53]
    two_complement_buffer_2_21 <= two_complement_2_21; // @[block_division.scala 216:53]
    two_complement_buffer_2_22 <= two_complement_2_22; // @[block_division.scala 216:53]
    two_complement_buffer_2_23 <= two_complement_2_23; // @[block_division.scala 216:53]
    two_complement_buffer_2_24 <= two_complement_2_24; // @[block_division.scala 216:53]
    two_complement_buffer_2_25 <= two_complement_2_25; // @[block_division.scala 216:53]
    two_complement_buffer_2_26 <= two_complement_2_26; // @[block_division.scala 216:53]
    two_complement_buffer_2_27 <= two_complement_2_27; // @[block_division.scala 216:53]
    two_complement_buffer_2_28 <= two_complement_2_28; // @[block_division.scala 216:53]
    two_complement_buffer_2_29 <= two_complement_2_29; // @[block_division.scala 216:53]
    two_complement_buffer_2_30 <= two_complement_2_30; // @[block_division.scala 216:53]
    two_complement_buffer_2_31 <= two_complement_2_31; // @[block_division.scala 216:53]
    two_complement_buffer_2_32 <= two_complement_2_32; // @[block_division.scala 216:53]
    two_complement_buffer_2_33 <= two_complement_2_33; // @[block_division.scala 216:53]
    two_complement_buffer_2_34 <= two_complement_2_34; // @[block_division.scala 216:53]
    two_complement_buffer_2_35 <= two_complement_2_35; // @[block_division.scala 216:53]
    two_complement_buffer_2_36 <= two_complement_2_36; // @[block_division.scala 216:53]
    two_complement_buffer_2_37 <= two_complement_2_37; // @[block_division.scala 216:53]
    two_complement_buffer_2_38 <= two_complement_2_38; // @[block_division.scala 216:53]
    two_complement_buffer_2_39 <= two_complement_2_39; // @[block_division.scala 216:53]
    two_complement_buffer_2_40 <= two_complement_2_40; // @[block_division.scala 216:53]
    two_complement_buffer_2_41 <= two_complement_2_41; // @[block_division.scala 216:53]
    two_complement_buffer_2_42 <= two_complement_2_42; // @[block_division.scala 216:53]
    two_complement_buffer_2_43 <= two_complement_2_43; // @[block_division.scala 216:53]
    two_complement_buffer_2_44 <= two_complement_2_44; // @[block_division.scala 216:53]
    two_complement_buffer_2_45 <= two_complement_2_45; // @[block_division.scala 216:53]
    two_complement_buffer_2_46 <= two_complement_2_46; // @[block_division.scala 216:53]
    two_complement_buffer_2_47 <= two_complement_2_47; // @[block_division.scala 216:53]
    two_complement_buffer_2_48 <= two_complement_2_48; // @[block_division.scala 216:53]
    two_complement_buffer_2_49 <= two_complement_2_49; // @[block_division.scala 216:53]
    two_complement_buffer_2_50 <= two_complement_2_50; // @[block_division.scala 216:53]
    two_complement_buffer_2_51 <= two_complement_2_51; // @[block_division.scala 216:53]
    two_complement_buffer_2_52 <= two_complement_2_52; // @[block_division.scala 216:53]
    two_complement_buffer_2_53 <= two_complement_2_53; // @[block_division.scala 216:53]
    two_complement_buffer_2_54 <= two_complement_2_54; // @[block_division.scala 216:53]
    two_complement_buffer_2_55 <= two_complement_2_55; // @[block_division.scala 216:53]
    two_complement_buffer_2_56 <= two_complement_2_56; // @[block_division.scala 216:53]
    two_complement_buffer_2_57 <= two_complement_2_57; // @[block_division.scala 216:53]
    two_complement_buffer_2_58 <= two_complement_2_58; // @[block_division.scala 216:53]
    two_complement_buffer_2_59 <= two_complement_2_59; // @[block_division.scala 216:53]
    two_complement_buffer_2_60 <= two_complement_2_60; // @[block_division.scala 216:53]
    two_complement_buffer_2_61 <= two_complement_2_61; // @[block_division.scala 216:53]
    two_complement_buffer_2_62 <= two_complement_2_62; // @[block_division.scala 216:53]
    two_complement_buffer_2_63 <= two_complement_2_63; // @[block_division.scala 216:53]
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_128 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_128 <= io_man_a_128; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_128 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_128 <= io_sign_a_128; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_129 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_129 <= io_man_a_129; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_129 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_129 <= io_sign_a_129; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_130 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_130 <= io_man_a_130; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_130 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_130 <= io_sign_a_130; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_131 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_131 <= io_man_a_131; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_131 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_131 <= io_sign_a_131; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_132 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_132 <= io_man_a_132; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_132 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_132 <= io_sign_a_132; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_133 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_133 <= io_man_a_133; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_133 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_133 <= io_sign_a_133; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_134 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_134 <= io_man_a_134; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_134 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_134 <= io_sign_a_134; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_135 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_135 <= io_man_a_135; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_135 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_135 <= io_sign_a_135; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_136 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_136 <= io_man_a_136; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_136 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_136 <= io_sign_a_136; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_137 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_137 <= io_man_a_137; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_137 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_137 <= io_sign_a_137; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_138 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_138 <= io_man_a_138; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_138 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_138 <= io_sign_a_138; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_139 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_139 <= io_man_a_139; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_139 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_139 <= io_sign_a_139; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_140 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_140 <= io_man_a_140; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_140 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_140 <= io_sign_a_140; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_141 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_141 <= io_man_a_141; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_141 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_141 <= io_sign_a_141; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_142 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_142 <= io_man_a_142; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_142 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_142 <= io_sign_a_142; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_143 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_143 <= io_man_a_143; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_143 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_143 <= io_sign_a_143; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_144 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_144 <= io_man_a_144; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_144 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_144 <= io_sign_a_144; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_145 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_145 <= io_man_a_145; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_145 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_145 <= io_sign_a_145; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_146 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_146 <= io_man_a_146; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_146 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_146 <= io_sign_a_146; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_147 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_147 <= io_man_a_147; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_147 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_147 <= io_sign_a_147; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_148 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_148 <= io_man_a_148; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_148 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_148 <= io_sign_a_148; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_149 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_149 <= io_man_a_149; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_149 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_149 <= io_sign_a_149; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_150 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_150 <= io_man_a_150; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_150 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_150 <= io_sign_a_150; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_151 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_151 <= io_man_a_151; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_151 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_151 <= io_sign_a_151; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_152 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_152 <= io_man_a_152; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_152 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_152 <= io_sign_a_152; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_153 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_153 <= io_man_a_153; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_153 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_153 <= io_sign_a_153; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_154 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_154 <= io_man_a_154; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_154 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_154 <= io_sign_a_154; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_155 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_155 <= io_man_a_155; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_155 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_155 <= io_sign_a_155; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_156 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_156 <= io_man_a_156; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_156 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_156 <= io_sign_a_156; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_157 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_157 <= io_man_a_157; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_157 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_157 <= io_sign_a_157; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_158 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_158 <= io_man_a_158; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_158 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_158 <= io_sign_a_158; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_159 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_159 <= io_man_a_159; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_159 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_159 <= io_sign_a_159; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_160 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_160 <= io_man_a_160; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_160 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_160 <= io_sign_a_160; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_161 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_161 <= io_man_a_161; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_161 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_161 <= io_sign_a_161; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_162 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_162 <= io_man_a_162; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_162 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_162 <= io_sign_a_162; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_163 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_163 <= io_man_a_163; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_163 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_163 <= io_sign_a_163; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_164 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_164 <= io_man_a_164; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_164 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_164 <= io_sign_a_164; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_165 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_165 <= io_man_a_165; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_165 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_165 <= io_sign_a_165; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_166 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_166 <= io_man_a_166; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_166 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_166 <= io_sign_a_166; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_167 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_167 <= io_man_a_167; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_167 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_167 <= io_sign_a_167; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_168 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_168 <= io_man_a_168; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_168 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_168 <= io_sign_a_168; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_169 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_169 <= io_man_a_169; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_169 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_169 <= io_sign_a_169; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_170 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_170 <= io_man_a_170; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_170 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_170 <= io_sign_a_170; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_171 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_171 <= io_man_a_171; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_171 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_171 <= io_sign_a_171; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_172 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_172 <= io_man_a_172; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_172 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_172 <= io_sign_a_172; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_173 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_173 <= io_man_a_173; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_173 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_173 <= io_sign_a_173; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_174 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_174 <= io_man_a_174; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_174 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_174 <= io_sign_a_174; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_175 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_175 <= io_man_a_175; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_175 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_175 <= io_sign_a_175; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_176 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_176 <= io_man_a_176; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_176 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_176 <= io_sign_a_176; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_177 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_177 <= io_man_a_177; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_177 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_177 <= io_sign_a_177; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_178 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_178 <= io_man_a_178; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_178 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_178 <= io_sign_a_178; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_179 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_179 <= io_man_a_179; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_179 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_179 <= io_sign_a_179; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_180 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_180 <= io_man_a_180; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_180 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_180 <= io_sign_a_180; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_181 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_181 <= io_man_a_181; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_181 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_181 <= io_sign_a_181; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_182 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_182 <= io_man_a_182; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_182 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_182 <= io_sign_a_182; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_183 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_183 <= io_man_a_183; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_183 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_183 <= io_sign_a_183; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_184 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_184 <= io_man_a_184; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_184 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_184 <= io_sign_a_184; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_185 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_185 <= io_man_a_185; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_185 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_185 <= io_sign_a_185; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_186 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_186 <= io_man_a_186; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_186 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_186 <= io_sign_a_186; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_187 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_187 <= io_man_a_187; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_187 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_187 <= io_sign_a_187; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_188 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_188 <= io_man_a_188; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_188 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_188 <= io_sign_a_188; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_189 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_189 <= io_man_a_189; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_189 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_189 <= io_sign_a_189; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_190 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_190 <= io_man_a_190; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_190 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_190 <= io_sign_a_190; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_191 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_191 <= io_man_a_191; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_191 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_191 <= io_sign_a_191; // @[block_division.scala 206:15]
    end
    dotProductRegs_3_0 <= _dotProductRegs_0_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_1 <= _dotProductRegs_1_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_2 <= _dotProductRegs_2_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_3 <= _dotProductRegs_3_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_4 <= _dotProductRegs_4_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_5 <= _dotProductRegs_5_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_6 <= _dotProductRegs_6_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_7 <= _dotProductRegs_7_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_8 <= _dotProductRegs_8_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_9 <= _dotProductRegs_9_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_10 <= _dotProductRegs_10_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_11 <= _dotProductRegs_11_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_12 <= _dotProductRegs_12_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_13 <= _dotProductRegs_13_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_14 <= _dotProductRegs_14_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_15 <= _dotProductRegs_15_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_16 <= _dotProductRegs_16_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_17 <= _dotProductRegs_17_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_18 <= _dotProductRegs_18_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_19 <= _dotProductRegs_19_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_20 <= _dotProductRegs_20_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_21 <= _dotProductRegs_21_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_22 <= _dotProductRegs_22_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_23 <= _dotProductRegs_23_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_24 <= _dotProductRegs_24_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_25 <= _dotProductRegs_25_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_26 <= _dotProductRegs_26_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_27 <= _dotProductRegs_27_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_28 <= _dotProductRegs_28_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_29 <= _dotProductRegs_29_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_30 <= _dotProductRegs_30_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_31 <= _dotProductRegs_31_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_32 <= _dotProductRegs_32_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_33 <= _dotProductRegs_33_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_34 <= _dotProductRegs_34_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_35 <= _dotProductRegs_35_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_36 <= _dotProductRegs_36_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_37 <= _dotProductRegs_37_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_38 <= _dotProductRegs_38_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_39 <= _dotProductRegs_39_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_40 <= _dotProductRegs_40_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_41 <= _dotProductRegs_41_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_42 <= _dotProductRegs_42_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_43 <= _dotProductRegs_43_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_44 <= _dotProductRegs_44_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_45 <= _dotProductRegs_45_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_46 <= _dotProductRegs_46_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_47 <= _dotProductRegs_47_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_48 <= _dotProductRegs_48_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_49 <= _dotProductRegs_49_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_50 <= _dotProductRegs_50_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_51 <= _dotProductRegs_51_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_52 <= _dotProductRegs_52_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_53 <= _dotProductRegs_53_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_54 <= _dotProductRegs_54_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_55 <= _dotProductRegs_55_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_56 <= _dotProductRegs_56_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_57 <= _dotProductRegs_57_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_58 <= _dotProductRegs_58_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_59 <= _dotProductRegs_59_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_60 <= _dotProductRegs_60_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_61 <= _dotProductRegs_61_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_62 <= _dotProductRegs_62_T_23[4:0]; // @[block_division.scala 209:25]
    dotProductRegs_3_63 <= _dotProductRegs_63_T_23[4:0]; // @[block_division.scala 209:25]
    signs_3_0 <= signReg_192 ^ io_sign_b_192; // @[block_division.scala 210:27]
    signs_3_1 <= signReg_193 ^ io_sign_b_193; // @[block_division.scala 210:27]
    signs_3_2 <= signReg_194 ^ io_sign_b_194; // @[block_division.scala 210:27]
    signs_3_3 <= signReg_195 ^ io_sign_b_195; // @[block_division.scala 210:27]
    signs_3_4 <= signReg_196 ^ io_sign_b_196; // @[block_division.scala 210:27]
    signs_3_5 <= signReg_197 ^ io_sign_b_197; // @[block_division.scala 210:27]
    signs_3_6 <= signReg_198 ^ io_sign_b_198; // @[block_division.scala 210:27]
    signs_3_7 <= signReg_199 ^ io_sign_b_199; // @[block_division.scala 210:27]
    signs_3_8 <= signReg_200 ^ io_sign_b_200; // @[block_division.scala 210:27]
    signs_3_9 <= signReg_201 ^ io_sign_b_201; // @[block_division.scala 210:27]
    signs_3_10 <= signReg_202 ^ io_sign_b_202; // @[block_division.scala 210:27]
    signs_3_11 <= signReg_203 ^ io_sign_b_203; // @[block_division.scala 210:27]
    signs_3_12 <= signReg_204 ^ io_sign_b_204; // @[block_division.scala 210:27]
    signs_3_13 <= signReg_205 ^ io_sign_b_205; // @[block_division.scala 210:27]
    signs_3_14 <= signReg_206 ^ io_sign_b_206; // @[block_division.scala 210:27]
    signs_3_15 <= signReg_207 ^ io_sign_b_207; // @[block_division.scala 210:27]
    signs_3_16 <= signReg_208 ^ io_sign_b_208; // @[block_division.scala 210:27]
    signs_3_17 <= signReg_209 ^ io_sign_b_209; // @[block_division.scala 210:27]
    signs_3_18 <= signReg_210 ^ io_sign_b_210; // @[block_division.scala 210:27]
    signs_3_19 <= signReg_211 ^ io_sign_b_211; // @[block_division.scala 210:27]
    signs_3_20 <= signReg_212 ^ io_sign_b_212; // @[block_division.scala 210:27]
    signs_3_21 <= signReg_213 ^ io_sign_b_213; // @[block_division.scala 210:27]
    signs_3_22 <= signReg_214 ^ io_sign_b_214; // @[block_division.scala 210:27]
    signs_3_23 <= signReg_215 ^ io_sign_b_215; // @[block_division.scala 210:27]
    signs_3_24 <= signReg_216 ^ io_sign_b_216; // @[block_division.scala 210:27]
    signs_3_25 <= signReg_217 ^ io_sign_b_217; // @[block_division.scala 210:27]
    signs_3_26 <= signReg_218 ^ io_sign_b_218; // @[block_division.scala 210:27]
    signs_3_27 <= signReg_219 ^ io_sign_b_219; // @[block_division.scala 210:27]
    signs_3_28 <= signReg_220 ^ io_sign_b_220; // @[block_division.scala 210:27]
    signs_3_29 <= signReg_221 ^ io_sign_b_221; // @[block_division.scala 210:27]
    signs_3_30 <= signReg_222 ^ io_sign_b_222; // @[block_division.scala 210:27]
    signs_3_31 <= signReg_223 ^ io_sign_b_223; // @[block_division.scala 210:27]
    signs_3_32 <= signReg_224 ^ io_sign_b_224; // @[block_division.scala 210:27]
    signs_3_33 <= signReg_225 ^ io_sign_b_225; // @[block_division.scala 210:27]
    signs_3_34 <= signReg_226 ^ io_sign_b_226; // @[block_division.scala 210:27]
    signs_3_35 <= signReg_227 ^ io_sign_b_227; // @[block_division.scala 210:27]
    signs_3_36 <= signReg_228 ^ io_sign_b_228; // @[block_division.scala 210:27]
    signs_3_37 <= signReg_229 ^ io_sign_b_229; // @[block_division.scala 210:27]
    signs_3_38 <= signReg_230 ^ io_sign_b_230; // @[block_division.scala 210:27]
    signs_3_39 <= signReg_231 ^ io_sign_b_231; // @[block_division.scala 210:27]
    signs_3_40 <= signReg_232 ^ io_sign_b_232; // @[block_division.scala 210:27]
    signs_3_41 <= signReg_233 ^ io_sign_b_233; // @[block_division.scala 210:27]
    signs_3_42 <= signReg_234 ^ io_sign_b_234; // @[block_division.scala 210:27]
    signs_3_43 <= signReg_235 ^ io_sign_b_235; // @[block_division.scala 210:27]
    signs_3_44 <= signReg_236 ^ io_sign_b_236; // @[block_division.scala 210:27]
    signs_3_45 <= signReg_237 ^ io_sign_b_237; // @[block_division.scala 210:27]
    signs_3_46 <= signReg_238 ^ io_sign_b_238; // @[block_division.scala 210:27]
    signs_3_47 <= signReg_239 ^ io_sign_b_239; // @[block_division.scala 210:27]
    signs_3_48 <= signReg_240 ^ io_sign_b_240; // @[block_division.scala 210:27]
    signs_3_49 <= signReg_241 ^ io_sign_b_241; // @[block_division.scala 210:27]
    signs_3_50 <= signReg_242 ^ io_sign_b_242; // @[block_division.scala 210:27]
    signs_3_51 <= signReg_243 ^ io_sign_b_243; // @[block_division.scala 210:27]
    signs_3_52 <= signReg_244 ^ io_sign_b_244; // @[block_division.scala 210:27]
    signs_3_53 <= signReg_245 ^ io_sign_b_245; // @[block_division.scala 210:27]
    signs_3_54 <= signReg_246 ^ io_sign_b_246; // @[block_division.scala 210:27]
    signs_3_55 <= signReg_247 ^ io_sign_b_247; // @[block_division.scala 210:27]
    signs_3_56 <= signReg_248 ^ io_sign_b_248; // @[block_division.scala 210:27]
    signs_3_57 <= signReg_249 ^ io_sign_b_249; // @[block_division.scala 210:27]
    signs_3_58 <= signReg_250 ^ io_sign_b_250; // @[block_division.scala 210:27]
    signs_3_59 <= signReg_251 ^ io_sign_b_251; // @[block_division.scala 210:27]
    signs_3_60 <= signReg_252 ^ io_sign_b_252; // @[block_division.scala 210:27]
    signs_3_61 <= signReg_253 ^ io_sign_b_253; // @[block_division.scala 210:27]
    signs_3_62 <= signReg_254 ^ io_sign_b_254; // @[block_division.scala 210:27]
    signs_3_63 <= signReg_255 ^ io_sign_b_255; // @[block_division.scala 210:27]
    if (signs_3_0) begin // @[block_division.scala 211:31]
      two_complement_3_0 <= _two_complement_0_T_25;
    end else begin
      two_complement_3_0 <= _two_complement_0_T_22;
    end
    if (signs_3_1) begin // @[block_division.scala 211:31]
      two_complement_3_1 <= _two_complement_1_T_25;
    end else begin
      two_complement_3_1 <= _two_complement_1_T_22;
    end
    if (signs_3_2) begin // @[block_division.scala 211:31]
      two_complement_3_2 <= _two_complement_2_T_25;
    end else begin
      two_complement_3_2 <= _two_complement_2_T_22;
    end
    if (signs_3_3) begin // @[block_division.scala 211:31]
      two_complement_3_3 <= _two_complement_3_T_25;
    end else begin
      two_complement_3_3 <= _two_complement_3_T_22;
    end
    if (signs_3_4) begin // @[block_division.scala 211:31]
      two_complement_3_4 <= _two_complement_4_T_25;
    end else begin
      two_complement_3_4 <= _two_complement_4_T_22;
    end
    if (signs_3_5) begin // @[block_division.scala 211:31]
      two_complement_3_5 <= _two_complement_5_T_25;
    end else begin
      two_complement_3_5 <= _two_complement_5_T_22;
    end
    if (signs_3_6) begin // @[block_division.scala 211:31]
      two_complement_3_6 <= _two_complement_6_T_25;
    end else begin
      two_complement_3_6 <= _two_complement_6_T_22;
    end
    if (signs_3_7) begin // @[block_division.scala 211:31]
      two_complement_3_7 <= _two_complement_7_T_25;
    end else begin
      two_complement_3_7 <= _two_complement_7_T_22;
    end
    if (signs_3_8) begin // @[block_division.scala 211:31]
      two_complement_3_8 <= _two_complement_8_T_25;
    end else begin
      two_complement_3_8 <= _two_complement_8_T_22;
    end
    if (signs_3_9) begin // @[block_division.scala 211:31]
      two_complement_3_9 <= _two_complement_9_T_25;
    end else begin
      two_complement_3_9 <= _two_complement_9_T_22;
    end
    if (signs_3_10) begin // @[block_division.scala 211:31]
      two_complement_3_10 <= _two_complement_10_T_25;
    end else begin
      two_complement_3_10 <= _two_complement_10_T_22;
    end
    if (signs_3_11) begin // @[block_division.scala 211:31]
      two_complement_3_11 <= _two_complement_11_T_25;
    end else begin
      two_complement_3_11 <= _two_complement_11_T_22;
    end
    if (signs_3_12) begin // @[block_division.scala 211:31]
      two_complement_3_12 <= _two_complement_12_T_25;
    end else begin
      two_complement_3_12 <= _two_complement_12_T_22;
    end
    if (signs_3_13) begin // @[block_division.scala 211:31]
      two_complement_3_13 <= _two_complement_13_T_25;
    end else begin
      two_complement_3_13 <= _two_complement_13_T_22;
    end
    if (signs_3_14) begin // @[block_division.scala 211:31]
      two_complement_3_14 <= _two_complement_14_T_25;
    end else begin
      two_complement_3_14 <= _two_complement_14_T_22;
    end
    if (signs_3_15) begin // @[block_division.scala 211:31]
      two_complement_3_15 <= _two_complement_15_T_25;
    end else begin
      two_complement_3_15 <= _two_complement_15_T_22;
    end
    if (signs_3_16) begin // @[block_division.scala 211:31]
      two_complement_3_16 <= _two_complement_16_T_25;
    end else begin
      two_complement_3_16 <= _two_complement_16_T_22;
    end
    if (signs_3_17) begin // @[block_division.scala 211:31]
      two_complement_3_17 <= _two_complement_17_T_25;
    end else begin
      two_complement_3_17 <= _two_complement_17_T_22;
    end
    if (signs_3_18) begin // @[block_division.scala 211:31]
      two_complement_3_18 <= _two_complement_18_T_25;
    end else begin
      two_complement_3_18 <= _two_complement_18_T_22;
    end
    if (signs_3_19) begin // @[block_division.scala 211:31]
      two_complement_3_19 <= _two_complement_19_T_25;
    end else begin
      two_complement_3_19 <= _two_complement_19_T_22;
    end
    if (signs_3_20) begin // @[block_division.scala 211:31]
      two_complement_3_20 <= _two_complement_20_T_25;
    end else begin
      two_complement_3_20 <= _two_complement_20_T_22;
    end
    if (signs_3_21) begin // @[block_division.scala 211:31]
      two_complement_3_21 <= _two_complement_21_T_25;
    end else begin
      two_complement_3_21 <= _two_complement_21_T_22;
    end
    if (signs_3_22) begin // @[block_division.scala 211:31]
      two_complement_3_22 <= _two_complement_22_T_25;
    end else begin
      two_complement_3_22 <= _two_complement_22_T_22;
    end
    if (signs_3_23) begin // @[block_division.scala 211:31]
      two_complement_3_23 <= _two_complement_23_T_25;
    end else begin
      two_complement_3_23 <= _two_complement_23_T_22;
    end
    if (signs_3_24) begin // @[block_division.scala 211:31]
      two_complement_3_24 <= _two_complement_24_T_25;
    end else begin
      two_complement_3_24 <= _two_complement_24_T_22;
    end
    if (signs_3_25) begin // @[block_division.scala 211:31]
      two_complement_3_25 <= _two_complement_25_T_25;
    end else begin
      two_complement_3_25 <= _two_complement_25_T_22;
    end
    if (signs_3_26) begin // @[block_division.scala 211:31]
      two_complement_3_26 <= _two_complement_26_T_25;
    end else begin
      two_complement_3_26 <= _two_complement_26_T_22;
    end
    if (signs_3_27) begin // @[block_division.scala 211:31]
      two_complement_3_27 <= _two_complement_27_T_25;
    end else begin
      two_complement_3_27 <= _two_complement_27_T_22;
    end
    if (signs_3_28) begin // @[block_division.scala 211:31]
      two_complement_3_28 <= _two_complement_28_T_25;
    end else begin
      two_complement_3_28 <= _two_complement_28_T_22;
    end
    if (signs_3_29) begin // @[block_division.scala 211:31]
      two_complement_3_29 <= _two_complement_29_T_25;
    end else begin
      two_complement_3_29 <= _two_complement_29_T_22;
    end
    if (signs_3_30) begin // @[block_division.scala 211:31]
      two_complement_3_30 <= _two_complement_30_T_25;
    end else begin
      two_complement_3_30 <= _two_complement_30_T_22;
    end
    if (signs_3_31) begin // @[block_division.scala 211:31]
      two_complement_3_31 <= _two_complement_31_T_25;
    end else begin
      two_complement_3_31 <= _two_complement_31_T_22;
    end
    if (signs_3_32) begin // @[block_division.scala 211:31]
      two_complement_3_32 <= _two_complement_32_T_25;
    end else begin
      two_complement_3_32 <= _two_complement_32_T_22;
    end
    if (signs_3_33) begin // @[block_division.scala 211:31]
      two_complement_3_33 <= _two_complement_33_T_25;
    end else begin
      two_complement_3_33 <= _two_complement_33_T_22;
    end
    if (signs_3_34) begin // @[block_division.scala 211:31]
      two_complement_3_34 <= _two_complement_34_T_25;
    end else begin
      two_complement_3_34 <= _two_complement_34_T_22;
    end
    if (signs_3_35) begin // @[block_division.scala 211:31]
      two_complement_3_35 <= _two_complement_35_T_25;
    end else begin
      two_complement_3_35 <= _two_complement_35_T_22;
    end
    if (signs_3_36) begin // @[block_division.scala 211:31]
      two_complement_3_36 <= _two_complement_36_T_25;
    end else begin
      two_complement_3_36 <= _two_complement_36_T_22;
    end
    if (signs_3_37) begin // @[block_division.scala 211:31]
      two_complement_3_37 <= _two_complement_37_T_25;
    end else begin
      two_complement_3_37 <= _two_complement_37_T_22;
    end
    if (signs_3_38) begin // @[block_division.scala 211:31]
      two_complement_3_38 <= _two_complement_38_T_25;
    end else begin
      two_complement_3_38 <= _two_complement_38_T_22;
    end
    if (signs_3_39) begin // @[block_division.scala 211:31]
      two_complement_3_39 <= _two_complement_39_T_25;
    end else begin
      two_complement_3_39 <= _two_complement_39_T_22;
    end
    if (signs_3_40) begin // @[block_division.scala 211:31]
      two_complement_3_40 <= _two_complement_40_T_25;
    end else begin
      two_complement_3_40 <= _two_complement_40_T_22;
    end
    if (signs_3_41) begin // @[block_division.scala 211:31]
      two_complement_3_41 <= _two_complement_41_T_25;
    end else begin
      two_complement_3_41 <= _two_complement_41_T_22;
    end
    if (signs_3_42) begin // @[block_division.scala 211:31]
      two_complement_3_42 <= _two_complement_42_T_25;
    end else begin
      two_complement_3_42 <= _two_complement_42_T_22;
    end
    if (signs_3_43) begin // @[block_division.scala 211:31]
      two_complement_3_43 <= _two_complement_43_T_25;
    end else begin
      two_complement_3_43 <= _two_complement_43_T_22;
    end
    if (signs_3_44) begin // @[block_division.scala 211:31]
      two_complement_3_44 <= _two_complement_44_T_25;
    end else begin
      two_complement_3_44 <= _two_complement_44_T_22;
    end
    if (signs_3_45) begin // @[block_division.scala 211:31]
      two_complement_3_45 <= _two_complement_45_T_25;
    end else begin
      two_complement_3_45 <= _two_complement_45_T_22;
    end
    if (signs_3_46) begin // @[block_division.scala 211:31]
      two_complement_3_46 <= _two_complement_46_T_25;
    end else begin
      two_complement_3_46 <= _two_complement_46_T_22;
    end
    if (signs_3_47) begin // @[block_division.scala 211:31]
      two_complement_3_47 <= _two_complement_47_T_25;
    end else begin
      two_complement_3_47 <= _two_complement_47_T_22;
    end
    if (signs_3_48) begin // @[block_division.scala 211:31]
      two_complement_3_48 <= _two_complement_48_T_25;
    end else begin
      two_complement_3_48 <= _two_complement_48_T_22;
    end
    if (signs_3_49) begin // @[block_division.scala 211:31]
      two_complement_3_49 <= _two_complement_49_T_25;
    end else begin
      two_complement_3_49 <= _two_complement_49_T_22;
    end
    if (signs_3_50) begin // @[block_division.scala 211:31]
      two_complement_3_50 <= _two_complement_50_T_25;
    end else begin
      two_complement_3_50 <= _two_complement_50_T_22;
    end
    if (signs_3_51) begin // @[block_division.scala 211:31]
      two_complement_3_51 <= _two_complement_51_T_25;
    end else begin
      two_complement_3_51 <= _two_complement_51_T_22;
    end
    if (signs_3_52) begin // @[block_division.scala 211:31]
      two_complement_3_52 <= _two_complement_52_T_25;
    end else begin
      two_complement_3_52 <= _two_complement_52_T_22;
    end
    if (signs_3_53) begin // @[block_division.scala 211:31]
      two_complement_3_53 <= _two_complement_53_T_25;
    end else begin
      two_complement_3_53 <= _two_complement_53_T_22;
    end
    if (signs_3_54) begin // @[block_division.scala 211:31]
      two_complement_3_54 <= _two_complement_54_T_25;
    end else begin
      two_complement_3_54 <= _two_complement_54_T_22;
    end
    if (signs_3_55) begin // @[block_division.scala 211:31]
      two_complement_3_55 <= _two_complement_55_T_25;
    end else begin
      two_complement_3_55 <= _two_complement_55_T_22;
    end
    if (signs_3_56) begin // @[block_division.scala 211:31]
      two_complement_3_56 <= _two_complement_56_T_25;
    end else begin
      two_complement_3_56 <= _two_complement_56_T_22;
    end
    if (signs_3_57) begin // @[block_division.scala 211:31]
      two_complement_3_57 <= _two_complement_57_T_25;
    end else begin
      two_complement_3_57 <= _two_complement_57_T_22;
    end
    if (signs_3_58) begin // @[block_division.scala 211:31]
      two_complement_3_58 <= _two_complement_58_T_25;
    end else begin
      two_complement_3_58 <= _two_complement_58_T_22;
    end
    if (signs_3_59) begin // @[block_division.scala 211:31]
      two_complement_3_59 <= _two_complement_59_T_25;
    end else begin
      two_complement_3_59 <= _two_complement_59_T_22;
    end
    if (signs_3_60) begin // @[block_division.scala 211:31]
      two_complement_3_60 <= _two_complement_60_T_25;
    end else begin
      two_complement_3_60 <= _two_complement_60_T_22;
    end
    if (signs_3_61) begin // @[block_division.scala 211:31]
      two_complement_3_61 <= _two_complement_61_T_25;
    end else begin
      two_complement_3_61 <= _two_complement_61_T_22;
    end
    if (signs_3_62) begin // @[block_division.scala 211:31]
      two_complement_3_62 <= _two_complement_62_T_25;
    end else begin
      two_complement_3_62 <= _two_complement_62_T_22;
    end
    if (signs_3_63) begin // @[block_division.scala 211:31]
      two_complement_3_63 <= _two_complement_63_T_25;
    end else begin
      two_complement_3_63 <= _two_complement_63_T_22;
    end
    two_complement_buffer_3_0 <= two_complement_3_0; // @[block_division.scala 216:53]
    two_complement_buffer_3_1 <= two_complement_3_1; // @[block_division.scala 216:53]
    two_complement_buffer_3_2 <= two_complement_3_2; // @[block_division.scala 216:53]
    two_complement_buffer_3_3 <= two_complement_3_3; // @[block_division.scala 216:53]
    two_complement_buffer_3_4 <= two_complement_3_4; // @[block_division.scala 216:53]
    two_complement_buffer_3_5 <= two_complement_3_5; // @[block_division.scala 216:53]
    two_complement_buffer_3_6 <= two_complement_3_6; // @[block_division.scala 216:53]
    two_complement_buffer_3_7 <= two_complement_3_7; // @[block_division.scala 216:53]
    two_complement_buffer_3_8 <= two_complement_3_8; // @[block_division.scala 216:53]
    two_complement_buffer_3_9 <= two_complement_3_9; // @[block_division.scala 216:53]
    two_complement_buffer_3_10 <= two_complement_3_10; // @[block_division.scala 216:53]
    two_complement_buffer_3_11 <= two_complement_3_11; // @[block_division.scala 216:53]
    two_complement_buffer_3_12 <= two_complement_3_12; // @[block_division.scala 216:53]
    two_complement_buffer_3_13 <= two_complement_3_13; // @[block_division.scala 216:53]
    two_complement_buffer_3_14 <= two_complement_3_14; // @[block_division.scala 216:53]
    two_complement_buffer_3_15 <= two_complement_3_15; // @[block_division.scala 216:53]
    two_complement_buffer_3_16 <= two_complement_3_16; // @[block_division.scala 216:53]
    two_complement_buffer_3_17 <= two_complement_3_17; // @[block_division.scala 216:53]
    two_complement_buffer_3_18 <= two_complement_3_18; // @[block_division.scala 216:53]
    two_complement_buffer_3_19 <= two_complement_3_19; // @[block_division.scala 216:53]
    two_complement_buffer_3_20 <= two_complement_3_20; // @[block_division.scala 216:53]
    two_complement_buffer_3_21 <= two_complement_3_21; // @[block_division.scala 216:53]
    two_complement_buffer_3_22 <= two_complement_3_22; // @[block_division.scala 216:53]
    two_complement_buffer_3_23 <= two_complement_3_23; // @[block_division.scala 216:53]
    two_complement_buffer_3_24 <= two_complement_3_24; // @[block_division.scala 216:53]
    two_complement_buffer_3_25 <= two_complement_3_25; // @[block_division.scala 216:53]
    two_complement_buffer_3_26 <= two_complement_3_26; // @[block_division.scala 216:53]
    two_complement_buffer_3_27 <= two_complement_3_27; // @[block_division.scala 216:53]
    two_complement_buffer_3_28 <= two_complement_3_28; // @[block_division.scala 216:53]
    two_complement_buffer_3_29 <= two_complement_3_29; // @[block_division.scala 216:53]
    two_complement_buffer_3_30 <= two_complement_3_30; // @[block_division.scala 216:53]
    two_complement_buffer_3_31 <= two_complement_3_31; // @[block_division.scala 216:53]
    two_complement_buffer_3_32 <= two_complement_3_32; // @[block_division.scala 216:53]
    two_complement_buffer_3_33 <= two_complement_3_33; // @[block_division.scala 216:53]
    two_complement_buffer_3_34 <= two_complement_3_34; // @[block_division.scala 216:53]
    two_complement_buffer_3_35 <= two_complement_3_35; // @[block_division.scala 216:53]
    two_complement_buffer_3_36 <= two_complement_3_36; // @[block_division.scala 216:53]
    two_complement_buffer_3_37 <= two_complement_3_37; // @[block_division.scala 216:53]
    two_complement_buffer_3_38 <= two_complement_3_38; // @[block_division.scala 216:53]
    two_complement_buffer_3_39 <= two_complement_3_39; // @[block_division.scala 216:53]
    two_complement_buffer_3_40 <= two_complement_3_40; // @[block_division.scala 216:53]
    two_complement_buffer_3_41 <= two_complement_3_41; // @[block_division.scala 216:53]
    two_complement_buffer_3_42 <= two_complement_3_42; // @[block_division.scala 216:53]
    two_complement_buffer_3_43 <= two_complement_3_43; // @[block_division.scala 216:53]
    two_complement_buffer_3_44 <= two_complement_3_44; // @[block_division.scala 216:53]
    two_complement_buffer_3_45 <= two_complement_3_45; // @[block_division.scala 216:53]
    two_complement_buffer_3_46 <= two_complement_3_46; // @[block_division.scala 216:53]
    two_complement_buffer_3_47 <= two_complement_3_47; // @[block_division.scala 216:53]
    two_complement_buffer_3_48 <= two_complement_3_48; // @[block_division.scala 216:53]
    two_complement_buffer_3_49 <= two_complement_3_49; // @[block_division.scala 216:53]
    two_complement_buffer_3_50 <= two_complement_3_50; // @[block_division.scala 216:53]
    two_complement_buffer_3_51 <= two_complement_3_51; // @[block_division.scala 216:53]
    two_complement_buffer_3_52 <= two_complement_3_52; // @[block_division.scala 216:53]
    two_complement_buffer_3_53 <= two_complement_3_53; // @[block_division.scala 216:53]
    two_complement_buffer_3_54 <= two_complement_3_54; // @[block_division.scala 216:53]
    two_complement_buffer_3_55 <= two_complement_3_55; // @[block_division.scala 216:53]
    two_complement_buffer_3_56 <= two_complement_3_56; // @[block_division.scala 216:53]
    two_complement_buffer_3_57 <= two_complement_3_57; // @[block_division.scala 216:53]
    two_complement_buffer_3_58 <= two_complement_3_58; // @[block_division.scala 216:53]
    two_complement_buffer_3_59 <= two_complement_3_59; // @[block_division.scala 216:53]
    two_complement_buffer_3_60 <= two_complement_3_60; // @[block_division.scala 216:53]
    two_complement_buffer_3_61 <= two_complement_3_61; // @[block_division.scala 216:53]
    two_complement_buffer_3_62 <= two_complement_3_62; // @[block_division.scala 216:53]
    two_complement_buffer_3_63 <= two_complement_3_63; // @[block_division.scala 216:53]
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_192 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_192 <= io_man_a_192; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_192 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_192 <= io_sign_a_192; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_193 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_193 <= io_man_a_193; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_193 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_193 <= io_sign_a_193; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_194 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_194 <= io_man_a_194; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_194 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_194 <= io_sign_a_194; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_195 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_195 <= io_man_a_195; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_195 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_195 <= io_sign_a_195; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_196 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_196 <= io_man_a_196; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_196 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_196 <= io_sign_a_196; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_197 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_197 <= io_man_a_197; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_197 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_197 <= io_sign_a_197; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_198 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_198 <= io_man_a_198; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_198 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_198 <= io_sign_a_198; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_199 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_199 <= io_man_a_199; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_199 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_199 <= io_sign_a_199; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_200 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_200 <= io_man_a_200; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_200 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_200 <= io_sign_a_200; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_201 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_201 <= io_man_a_201; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_201 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_201 <= io_sign_a_201; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_202 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_202 <= io_man_a_202; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_202 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_202 <= io_sign_a_202; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_203 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_203 <= io_man_a_203; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_203 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_203 <= io_sign_a_203; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_204 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_204 <= io_man_a_204; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_204 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_204 <= io_sign_a_204; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_205 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_205 <= io_man_a_205; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_205 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_205 <= io_sign_a_205; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_206 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_206 <= io_man_a_206; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_206 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_206 <= io_sign_a_206; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_207 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_207 <= io_man_a_207; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_207 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_207 <= io_sign_a_207; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_208 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_208 <= io_man_a_208; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_208 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_208 <= io_sign_a_208; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_209 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_209 <= io_man_a_209; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_209 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_209 <= io_sign_a_209; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_210 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_210 <= io_man_a_210; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_210 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_210 <= io_sign_a_210; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_211 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_211 <= io_man_a_211; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_211 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_211 <= io_sign_a_211; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_212 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_212 <= io_man_a_212; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_212 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_212 <= io_sign_a_212; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_213 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_213 <= io_man_a_213; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_213 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_213 <= io_sign_a_213; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_214 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_214 <= io_man_a_214; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_214 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_214 <= io_sign_a_214; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_215 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_215 <= io_man_a_215; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_215 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_215 <= io_sign_a_215; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_216 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_216 <= io_man_a_216; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_216 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_216 <= io_sign_a_216; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_217 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_217 <= io_man_a_217; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_217 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_217 <= io_sign_a_217; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_218 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_218 <= io_man_a_218; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_218 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_218 <= io_sign_a_218; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_219 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_219 <= io_man_a_219; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_219 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_219 <= io_sign_a_219; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_220 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_220 <= io_man_a_220; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_220 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_220 <= io_sign_a_220; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_221 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_221 <= io_man_a_221; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_221 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_221 <= io_sign_a_221; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_222 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_222 <= io_man_a_222; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_222 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_222 <= io_sign_a_222; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_223 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_223 <= io_man_a_223; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_223 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_223 <= io_sign_a_223; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_224 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_224 <= io_man_a_224; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_224 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_224 <= io_sign_a_224; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_225 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_225 <= io_man_a_225; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_225 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_225 <= io_sign_a_225; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_226 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_226 <= io_man_a_226; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_226 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_226 <= io_sign_a_226; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_227 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_227 <= io_man_a_227; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_227 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_227 <= io_sign_a_227; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_228 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_228 <= io_man_a_228; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_228 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_228 <= io_sign_a_228; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_229 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_229 <= io_man_a_229; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_229 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_229 <= io_sign_a_229; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_230 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_230 <= io_man_a_230; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_230 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_230 <= io_sign_a_230; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_231 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_231 <= io_man_a_231; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_231 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_231 <= io_sign_a_231; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_232 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_232 <= io_man_a_232; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_232 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_232 <= io_sign_a_232; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_233 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_233 <= io_man_a_233; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_233 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_233 <= io_sign_a_233; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_234 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_234 <= io_man_a_234; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_234 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_234 <= io_sign_a_234; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_235 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_235 <= io_man_a_235; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_235 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_235 <= io_sign_a_235; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_236 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_236 <= io_man_a_236; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_236 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_236 <= io_sign_a_236; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_237 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_237 <= io_man_a_237; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_237 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_237 <= io_sign_a_237; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_238 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_238 <= io_man_a_238; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_238 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_238 <= io_sign_a_238; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_239 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_239 <= io_man_a_239; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_239 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_239 <= io_sign_a_239; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_240 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_240 <= io_man_a_240; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_240 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_240 <= io_sign_a_240; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_241 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_241 <= io_man_a_241; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_241 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_241 <= io_sign_a_241; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_242 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_242 <= io_man_a_242; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_242 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_242 <= io_sign_a_242; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_243 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_243 <= io_man_a_243; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_243 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_243 <= io_sign_a_243; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_244 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_244 <= io_man_a_244; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_244 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_244 <= io_sign_a_244; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_245 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_245 <= io_man_a_245; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_245 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_245 <= io_sign_a_245; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_246 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_246 <= io_man_a_246; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_246 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_246 <= io_sign_a_246; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_247 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_247 <= io_man_a_247; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_247 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_247 <= io_sign_a_247; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_248 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_248 <= io_man_a_248; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_248 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_248 <= io_sign_a_248; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_249 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_249 <= io_man_a_249; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_249 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_249 <= io_sign_a_249; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_250 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_250 <= io_man_a_250; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_250 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_250 <= io_sign_a_250; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_251 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_251 <= io_man_a_251; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_251 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_251 <= io_sign_a_251; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_252 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_252 <= io_man_a_252; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_252 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_252 <= io_sign_a_252; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_253 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_253 <= io_man_a_253; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_253 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_253 <= io_sign_a_253; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_254 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_254 <= io_man_a_254; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_254 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_254 <= io_sign_a_254; // @[block_division.scala 206:15]
    end
    if (reset) begin // @[block_division.scala 204:34]
      multiplierReg_255 <= 5'h0; // @[block_division.scala 204:34]
    end else begin
      multiplierReg_255 <= io_man_a_255; // @[block_division.scala 207:21]
    end
    if (reset) begin // @[block_division.scala 205:28]
      signReg_255 <= 1'h0; // @[block_division.scala 205:28]
    end else begin
      signReg_255 <= io_sign_a_255; // @[block_division.scala 206:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  exp_output_0 = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  exp_output_1 = _RAND_1[8:0];
  _RAND_2 = {1{`RANDOM}};
  exp_output_2 = _RAND_2[8:0];
  _RAND_3 = {1{`RANDOM}};
  exp_output_3 = _RAND_3[8:0];
  _RAND_4 = {1{`RANDOM}};
  acc_0 = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  acc_1 = _RAND_5[5:0];
  _RAND_6 = {1{`RANDOM}};
  acc_2 = _RAND_6[5:0];
  _RAND_7 = {1{`RANDOM}};
  acc_3 = _RAND_7[5:0];
  _RAND_8 = {1{`RANDOM}};
  dotProductRegs__0 = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  dotProductRegs__1 = _RAND_9[4:0];
  _RAND_10 = {1{`RANDOM}};
  dotProductRegs__2 = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  dotProductRegs__3 = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  dotProductRegs__4 = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  dotProductRegs__5 = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  dotProductRegs__6 = _RAND_14[4:0];
  _RAND_15 = {1{`RANDOM}};
  dotProductRegs__7 = _RAND_15[4:0];
  _RAND_16 = {1{`RANDOM}};
  dotProductRegs__8 = _RAND_16[4:0];
  _RAND_17 = {1{`RANDOM}};
  dotProductRegs__9 = _RAND_17[4:0];
  _RAND_18 = {1{`RANDOM}};
  dotProductRegs__10 = _RAND_18[4:0];
  _RAND_19 = {1{`RANDOM}};
  dotProductRegs__11 = _RAND_19[4:0];
  _RAND_20 = {1{`RANDOM}};
  dotProductRegs__12 = _RAND_20[4:0];
  _RAND_21 = {1{`RANDOM}};
  dotProductRegs__13 = _RAND_21[4:0];
  _RAND_22 = {1{`RANDOM}};
  dotProductRegs__14 = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  dotProductRegs__15 = _RAND_23[4:0];
  _RAND_24 = {1{`RANDOM}};
  dotProductRegs__16 = _RAND_24[4:0];
  _RAND_25 = {1{`RANDOM}};
  dotProductRegs__17 = _RAND_25[4:0];
  _RAND_26 = {1{`RANDOM}};
  dotProductRegs__18 = _RAND_26[4:0];
  _RAND_27 = {1{`RANDOM}};
  dotProductRegs__19 = _RAND_27[4:0];
  _RAND_28 = {1{`RANDOM}};
  dotProductRegs__20 = _RAND_28[4:0];
  _RAND_29 = {1{`RANDOM}};
  dotProductRegs__21 = _RAND_29[4:0];
  _RAND_30 = {1{`RANDOM}};
  dotProductRegs__22 = _RAND_30[4:0];
  _RAND_31 = {1{`RANDOM}};
  dotProductRegs__23 = _RAND_31[4:0];
  _RAND_32 = {1{`RANDOM}};
  dotProductRegs__24 = _RAND_32[4:0];
  _RAND_33 = {1{`RANDOM}};
  dotProductRegs__25 = _RAND_33[4:0];
  _RAND_34 = {1{`RANDOM}};
  dotProductRegs__26 = _RAND_34[4:0];
  _RAND_35 = {1{`RANDOM}};
  dotProductRegs__27 = _RAND_35[4:0];
  _RAND_36 = {1{`RANDOM}};
  dotProductRegs__28 = _RAND_36[4:0];
  _RAND_37 = {1{`RANDOM}};
  dotProductRegs__29 = _RAND_37[4:0];
  _RAND_38 = {1{`RANDOM}};
  dotProductRegs__30 = _RAND_38[4:0];
  _RAND_39 = {1{`RANDOM}};
  dotProductRegs__31 = _RAND_39[4:0];
  _RAND_40 = {1{`RANDOM}};
  dotProductRegs__32 = _RAND_40[4:0];
  _RAND_41 = {1{`RANDOM}};
  dotProductRegs__33 = _RAND_41[4:0];
  _RAND_42 = {1{`RANDOM}};
  dotProductRegs__34 = _RAND_42[4:0];
  _RAND_43 = {1{`RANDOM}};
  dotProductRegs__35 = _RAND_43[4:0];
  _RAND_44 = {1{`RANDOM}};
  dotProductRegs__36 = _RAND_44[4:0];
  _RAND_45 = {1{`RANDOM}};
  dotProductRegs__37 = _RAND_45[4:0];
  _RAND_46 = {1{`RANDOM}};
  dotProductRegs__38 = _RAND_46[4:0];
  _RAND_47 = {1{`RANDOM}};
  dotProductRegs__39 = _RAND_47[4:0];
  _RAND_48 = {1{`RANDOM}};
  dotProductRegs__40 = _RAND_48[4:0];
  _RAND_49 = {1{`RANDOM}};
  dotProductRegs__41 = _RAND_49[4:0];
  _RAND_50 = {1{`RANDOM}};
  dotProductRegs__42 = _RAND_50[4:0];
  _RAND_51 = {1{`RANDOM}};
  dotProductRegs__43 = _RAND_51[4:0];
  _RAND_52 = {1{`RANDOM}};
  dotProductRegs__44 = _RAND_52[4:0];
  _RAND_53 = {1{`RANDOM}};
  dotProductRegs__45 = _RAND_53[4:0];
  _RAND_54 = {1{`RANDOM}};
  dotProductRegs__46 = _RAND_54[4:0];
  _RAND_55 = {1{`RANDOM}};
  dotProductRegs__47 = _RAND_55[4:0];
  _RAND_56 = {1{`RANDOM}};
  dotProductRegs__48 = _RAND_56[4:0];
  _RAND_57 = {1{`RANDOM}};
  dotProductRegs__49 = _RAND_57[4:0];
  _RAND_58 = {1{`RANDOM}};
  dotProductRegs__50 = _RAND_58[4:0];
  _RAND_59 = {1{`RANDOM}};
  dotProductRegs__51 = _RAND_59[4:0];
  _RAND_60 = {1{`RANDOM}};
  dotProductRegs__52 = _RAND_60[4:0];
  _RAND_61 = {1{`RANDOM}};
  dotProductRegs__53 = _RAND_61[4:0];
  _RAND_62 = {1{`RANDOM}};
  dotProductRegs__54 = _RAND_62[4:0];
  _RAND_63 = {1{`RANDOM}};
  dotProductRegs__55 = _RAND_63[4:0];
  _RAND_64 = {1{`RANDOM}};
  dotProductRegs__56 = _RAND_64[4:0];
  _RAND_65 = {1{`RANDOM}};
  dotProductRegs__57 = _RAND_65[4:0];
  _RAND_66 = {1{`RANDOM}};
  dotProductRegs__58 = _RAND_66[4:0];
  _RAND_67 = {1{`RANDOM}};
  dotProductRegs__59 = _RAND_67[4:0];
  _RAND_68 = {1{`RANDOM}};
  dotProductRegs__60 = _RAND_68[4:0];
  _RAND_69 = {1{`RANDOM}};
  dotProductRegs__61 = _RAND_69[4:0];
  _RAND_70 = {1{`RANDOM}};
  dotProductRegs__62 = _RAND_70[4:0];
  _RAND_71 = {1{`RANDOM}};
  dotProductRegs__63 = _RAND_71[4:0];
  _RAND_72 = {1{`RANDOM}};
  signs__0 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  signs__1 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  signs__2 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  signs__3 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  signs__4 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  signs__5 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  signs__6 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  signs__7 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  signs__8 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  signs__9 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  signs__10 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  signs__11 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  signs__12 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  signs__13 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  signs__14 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  signs__15 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  signs__16 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  signs__17 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  signs__18 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  signs__19 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  signs__20 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  signs__21 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  signs__22 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  signs__23 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  signs__24 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  signs__25 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  signs__26 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  signs__27 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  signs__28 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  signs__29 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  signs__30 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  signs__31 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  signs__32 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  signs__33 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  signs__34 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  signs__35 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  signs__36 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  signs__37 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  signs__38 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  signs__39 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  signs__40 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  signs__41 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  signs__42 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  signs__43 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  signs__44 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  signs__45 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  signs__46 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  signs__47 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  signs__48 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  signs__49 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  signs__50 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  signs__51 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  signs__52 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  signs__53 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  signs__54 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  signs__55 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  signs__56 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  signs__57 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  signs__58 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  signs__59 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  signs__60 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  signs__61 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  signs__62 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  signs__63 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  two_complement__0 = _RAND_136[5:0];
  _RAND_137 = {1{`RANDOM}};
  two_complement__1 = _RAND_137[5:0];
  _RAND_138 = {1{`RANDOM}};
  two_complement__2 = _RAND_138[5:0];
  _RAND_139 = {1{`RANDOM}};
  two_complement__3 = _RAND_139[5:0];
  _RAND_140 = {1{`RANDOM}};
  two_complement__4 = _RAND_140[5:0];
  _RAND_141 = {1{`RANDOM}};
  two_complement__5 = _RAND_141[5:0];
  _RAND_142 = {1{`RANDOM}};
  two_complement__6 = _RAND_142[5:0];
  _RAND_143 = {1{`RANDOM}};
  two_complement__7 = _RAND_143[5:0];
  _RAND_144 = {1{`RANDOM}};
  two_complement__8 = _RAND_144[5:0];
  _RAND_145 = {1{`RANDOM}};
  two_complement__9 = _RAND_145[5:0];
  _RAND_146 = {1{`RANDOM}};
  two_complement__10 = _RAND_146[5:0];
  _RAND_147 = {1{`RANDOM}};
  two_complement__11 = _RAND_147[5:0];
  _RAND_148 = {1{`RANDOM}};
  two_complement__12 = _RAND_148[5:0];
  _RAND_149 = {1{`RANDOM}};
  two_complement__13 = _RAND_149[5:0];
  _RAND_150 = {1{`RANDOM}};
  two_complement__14 = _RAND_150[5:0];
  _RAND_151 = {1{`RANDOM}};
  two_complement__15 = _RAND_151[5:0];
  _RAND_152 = {1{`RANDOM}};
  two_complement__16 = _RAND_152[5:0];
  _RAND_153 = {1{`RANDOM}};
  two_complement__17 = _RAND_153[5:0];
  _RAND_154 = {1{`RANDOM}};
  two_complement__18 = _RAND_154[5:0];
  _RAND_155 = {1{`RANDOM}};
  two_complement__19 = _RAND_155[5:0];
  _RAND_156 = {1{`RANDOM}};
  two_complement__20 = _RAND_156[5:0];
  _RAND_157 = {1{`RANDOM}};
  two_complement__21 = _RAND_157[5:0];
  _RAND_158 = {1{`RANDOM}};
  two_complement__22 = _RAND_158[5:0];
  _RAND_159 = {1{`RANDOM}};
  two_complement__23 = _RAND_159[5:0];
  _RAND_160 = {1{`RANDOM}};
  two_complement__24 = _RAND_160[5:0];
  _RAND_161 = {1{`RANDOM}};
  two_complement__25 = _RAND_161[5:0];
  _RAND_162 = {1{`RANDOM}};
  two_complement__26 = _RAND_162[5:0];
  _RAND_163 = {1{`RANDOM}};
  two_complement__27 = _RAND_163[5:0];
  _RAND_164 = {1{`RANDOM}};
  two_complement__28 = _RAND_164[5:0];
  _RAND_165 = {1{`RANDOM}};
  two_complement__29 = _RAND_165[5:0];
  _RAND_166 = {1{`RANDOM}};
  two_complement__30 = _RAND_166[5:0];
  _RAND_167 = {1{`RANDOM}};
  two_complement__31 = _RAND_167[5:0];
  _RAND_168 = {1{`RANDOM}};
  two_complement__32 = _RAND_168[5:0];
  _RAND_169 = {1{`RANDOM}};
  two_complement__33 = _RAND_169[5:0];
  _RAND_170 = {1{`RANDOM}};
  two_complement__34 = _RAND_170[5:0];
  _RAND_171 = {1{`RANDOM}};
  two_complement__35 = _RAND_171[5:0];
  _RAND_172 = {1{`RANDOM}};
  two_complement__36 = _RAND_172[5:0];
  _RAND_173 = {1{`RANDOM}};
  two_complement__37 = _RAND_173[5:0];
  _RAND_174 = {1{`RANDOM}};
  two_complement__38 = _RAND_174[5:0];
  _RAND_175 = {1{`RANDOM}};
  two_complement__39 = _RAND_175[5:0];
  _RAND_176 = {1{`RANDOM}};
  two_complement__40 = _RAND_176[5:0];
  _RAND_177 = {1{`RANDOM}};
  two_complement__41 = _RAND_177[5:0];
  _RAND_178 = {1{`RANDOM}};
  two_complement__42 = _RAND_178[5:0];
  _RAND_179 = {1{`RANDOM}};
  two_complement__43 = _RAND_179[5:0];
  _RAND_180 = {1{`RANDOM}};
  two_complement__44 = _RAND_180[5:0];
  _RAND_181 = {1{`RANDOM}};
  two_complement__45 = _RAND_181[5:0];
  _RAND_182 = {1{`RANDOM}};
  two_complement__46 = _RAND_182[5:0];
  _RAND_183 = {1{`RANDOM}};
  two_complement__47 = _RAND_183[5:0];
  _RAND_184 = {1{`RANDOM}};
  two_complement__48 = _RAND_184[5:0];
  _RAND_185 = {1{`RANDOM}};
  two_complement__49 = _RAND_185[5:0];
  _RAND_186 = {1{`RANDOM}};
  two_complement__50 = _RAND_186[5:0];
  _RAND_187 = {1{`RANDOM}};
  two_complement__51 = _RAND_187[5:0];
  _RAND_188 = {1{`RANDOM}};
  two_complement__52 = _RAND_188[5:0];
  _RAND_189 = {1{`RANDOM}};
  two_complement__53 = _RAND_189[5:0];
  _RAND_190 = {1{`RANDOM}};
  two_complement__54 = _RAND_190[5:0];
  _RAND_191 = {1{`RANDOM}};
  two_complement__55 = _RAND_191[5:0];
  _RAND_192 = {1{`RANDOM}};
  two_complement__56 = _RAND_192[5:0];
  _RAND_193 = {1{`RANDOM}};
  two_complement__57 = _RAND_193[5:0];
  _RAND_194 = {1{`RANDOM}};
  two_complement__58 = _RAND_194[5:0];
  _RAND_195 = {1{`RANDOM}};
  two_complement__59 = _RAND_195[5:0];
  _RAND_196 = {1{`RANDOM}};
  two_complement__60 = _RAND_196[5:0];
  _RAND_197 = {1{`RANDOM}};
  two_complement__61 = _RAND_197[5:0];
  _RAND_198 = {1{`RANDOM}};
  two_complement__62 = _RAND_198[5:0];
  _RAND_199 = {1{`RANDOM}};
  two_complement__63 = _RAND_199[5:0];
  _RAND_200 = {1{`RANDOM}};
  two_complement_buffer__0 = _RAND_200[5:0];
  _RAND_201 = {1{`RANDOM}};
  two_complement_buffer__1 = _RAND_201[5:0];
  _RAND_202 = {1{`RANDOM}};
  two_complement_buffer__2 = _RAND_202[5:0];
  _RAND_203 = {1{`RANDOM}};
  two_complement_buffer__3 = _RAND_203[5:0];
  _RAND_204 = {1{`RANDOM}};
  two_complement_buffer__4 = _RAND_204[5:0];
  _RAND_205 = {1{`RANDOM}};
  two_complement_buffer__5 = _RAND_205[5:0];
  _RAND_206 = {1{`RANDOM}};
  two_complement_buffer__6 = _RAND_206[5:0];
  _RAND_207 = {1{`RANDOM}};
  two_complement_buffer__7 = _RAND_207[5:0];
  _RAND_208 = {1{`RANDOM}};
  two_complement_buffer__8 = _RAND_208[5:0];
  _RAND_209 = {1{`RANDOM}};
  two_complement_buffer__9 = _RAND_209[5:0];
  _RAND_210 = {1{`RANDOM}};
  two_complement_buffer__10 = _RAND_210[5:0];
  _RAND_211 = {1{`RANDOM}};
  two_complement_buffer__11 = _RAND_211[5:0];
  _RAND_212 = {1{`RANDOM}};
  two_complement_buffer__12 = _RAND_212[5:0];
  _RAND_213 = {1{`RANDOM}};
  two_complement_buffer__13 = _RAND_213[5:0];
  _RAND_214 = {1{`RANDOM}};
  two_complement_buffer__14 = _RAND_214[5:0];
  _RAND_215 = {1{`RANDOM}};
  two_complement_buffer__15 = _RAND_215[5:0];
  _RAND_216 = {1{`RANDOM}};
  two_complement_buffer__16 = _RAND_216[5:0];
  _RAND_217 = {1{`RANDOM}};
  two_complement_buffer__17 = _RAND_217[5:0];
  _RAND_218 = {1{`RANDOM}};
  two_complement_buffer__18 = _RAND_218[5:0];
  _RAND_219 = {1{`RANDOM}};
  two_complement_buffer__19 = _RAND_219[5:0];
  _RAND_220 = {1{`RANDOM}};
  two_complement_buffer__20 = _RAND_220[5:0];
  _RAND_221 = {1{`RANDOM}};
  two_complement_buffer__21 = _RAND_221[5:0];
  _RAND_222 = {1{`RANDOM}};
  two_complement_buffer__22 = _RAND_222[5:0];
  _RAND_223 = {1{`RANDOM}};
  two_complement_buffer__23 = _RAND_223[5:0];
  _RAND_224 = {1{`RANDOM}};
  two_complement_buffer__24 = _RAND_224[5:0];
  _RAND_225 = {1{`RANDOM}};
  two_complement_buffer__25 = _RAND_225[5:0];
  _RAND_226 = {1{`RANDOM}};
  two_complement_buffer__26 = _RAND_226[5:0];
  _RAND_227 = {1{`RANDOM}};
  two_complement_buffer__27 = _RAND_227[5:0];
  _RAND_228 = {1{`RANDOM}};
  two_complement_buffer__28 = _RAND_228[5:0];
  _RAND_229 = {1{`RANDOM}};
  two_complement_buffer__29 = _RAND_229[5:0];
  _RAND_230 = {1{`RANDOM}};
  two_complement_buffer__30 = _RAND_230[5:0];
  _RAND_231 = {1{`RANDOM}};
  two_complement_buffer__31 = _RAND_231[5:0];
  _RAND_232 = {1{`RANDOM}};
  two_complement_buffer__32 = _RAND_232[5:0];
  _RAND_233 = {1{`RANDOM}};
  two_complement_buffer__33 = _RAND_233[5:0];
  _RAND_234 = {1{`RANDOM}};
  two_complement_buffer__34 = _RAND_234[5:0];
  _RAND_235 = {1{`RANDOM}};
  two_complement_buffer__35 = _RAND_235[5:0];
  _RAND_236 = {1{`RANDOM}};
  two_complement_buffer__36 = _RAND_236[5:0];
  _RAND_237 = {1{`RANDOM}};
  two_complement_buffer__37 = _RAND_237[5:0];
  _RAND_238 = {1{`RANDOM}};
  two_complement_buffer__38 = _RAND_238[5:0];
  _RAND_239 = {1{`RANDOM}};
  two_complement_buffer__39 = _RAND_239[5:0];
  _RAND_240 = {1{`RANDOM}};
  two_complement_buffer__40 = _RAND_240[5:0];
  _RAND_241 = {1{`RANDOM}};
  two_complement_buffer__41 = _RAND_241[5:0];
  _RAND_242 = {1{`RANDOM}};
  two_complement_buffer__42 = _RAND_242[5:0];
  _RAND_243 = {1{`RANDOM}};
  two_complement_buffer__43 = _RAND_243[5:0];
  _RAND_244 = {1{`RANDOM}};
  two_complement_buffer__44 = _RAND_244[5:0];
  _RAND_245 = {1{`RANDOM}};
  two_complement_buffer__45 = _RAND_245[5:0];
  _RAND_246 = {1{`RANDOM}};
  two_complement_buffer__46 = _RAND_246[5:0];
  _RAND_247 = {1{`RANDOM}};
  two_complement_buffer__47 = _RAND_247[5:0];
  _RAND_248 = {1{`RANDOM}};
  two_complement_buffer__48 = _RAND_248[5:0];
  _RAND_249 = {1{`RANDOM}};
  two_complement_buffer__49 = _RAND_249[5:0];
  _RAND_250 = {1{`RANDOM}};
  two_complement_buffer__50 = _RAND_250[5:0];
  _RAND_251 = {1{`RANDOM}};
  two_complement_buffer__51 = _RAND_251[5:0];
  _RAND_252 = {1{`RANDOM}};
  two_complement_buffer__52 = _RAND_252[5:0];
  _RAND_253 = {1{`RANDOM}};
  two_complement_buffer__53 = _RAND_253[5:0];
  _RAND_254 = {1{`RANDOM}};
  two_complement_buffer__54 = _RAND_254[5:0];
  _RAND_255 = {1{`RANDOM}};
  two_complement_buffer__55 = _RAND_255[5:0];
  _RAND_256 = {1{`RANDOM}};
  two_complement_buffer__56 = _RAND_256[5:0];
  _RAND_257 = {1{`RANDOM}};
  two_complement_buffer__57 = _RAND_257[5:0];
  _RAND_258 = {1{`RANDOM}};
  two_complement_buffer__58 = _RAND_258[5:0];
  _RAND_259 = {1{`RANDOM}};
  two_complement_buffer__59 = _RAND_259[5:0];
  _RAND_260 = {1{`RANDOM}};
  two_complement_buffer__60 = _RAND_260[5:0];
  _RAND_261 = {1{`RANDOM}};
  two_complement_buffer__61 = _RAND_261[5:0];
  _RAND_262 = {1{`RANDOM}};
  two_complement_buffer__62 = _RAND_262[5:0];
  _RAND_263 = {1{`RANDOM}};
  two_complement_buffer__63 = _RAND_263[5:0];
  _RAND_264 = {1{`RANDOM}};
  multiplierReg = _RAND_264[4:0];
  _RAND_265 = {1{`RANDOM}};
  signReg = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  multiplierReg_1 = _RAND_266[4:0];
  _RAND_267 = {1{`RANDOM}};
  signReg_1 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  multiplierReg_2 = _RAND_268[4:0];
  _RAND_269 = {1{`RANDOM}};
  signReg_2 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  multiplierReg_3 = _RAND_270[4:0];
  _RAND_271 = {1{`RANDOM}};
  signReg_3 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  multiplierReg_4 = _RAND_272[4:0];
  _RAND_273 = {1{`RANDOM}};
  signReg_4 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  multiplierReg_5 = _RAND_274[4:0];
  _RAND_275 = {1{`RANDOM}};
  signReg_5 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  multiplierReg_6 = _RAND_276[4:0];
  _RAND_277 = {1{`RANDOM}};
  signReg_6 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  multiplierReg_7 = _RAND_278[4:0];
  _RAND_279 = {1{`RANDOM}};
  signReg_7 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  multiplierReg_8 = _RAND_280[4:0];
  _RAND_281 = {1{`RANDOM}};
  signReg_8 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  multiplierReg_9 = _RAND_282[4:0];
  _RAND_283 = {1{`RANDOM}};
  signReg_9 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  multiplierReg_10 = _RAND_284[4:0];
  _RAND_285 = {1{`RANDOM}};
  signReg_10 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  multiplierReg_11 = _RAND_286[4:0];
  _RAND_287 = {1{`RANDOM}};
  signReg_11 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  multiplierReg_12 = _RAND_288[4:0];
  _RAND_289 = {1{`RANDOM}};
  signReg_12 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  multiplierReg_13 = _RAND_290[4:0];
  _RAND_291 = {1{`RANDOM}};
  signReg_13 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  multiplierReg_14 = _RAND_292[4:0];
  _RAND_293 = {1{`RANDOM}};
  signReg_14 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  multiplierReg_15 = _RAND_294[4:0];
  _RAND_295 = {1{`RANDOM}};
  signReg_15 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  multiplierReg_16 = _RAND_296[4:0];
  _RAND_297 = {1{`RANDOM}};
  signReg_16 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  multiplierReg_17 = _RAND_298[4:0];
  _RAND_299 = {1{`RANDOM}};
  signReg_17 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  multiplierReg_18 = _RAND_300[4:0];
  _RAND_301 = {1{`RANDOM}};
  signReg_18 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  multiplierReg_19 = _RAND_302[4:0];
  _RAND_303 = {1{`RANDOM}};
  signReg_19 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  multiplierReg_20 = _RAND_304[4:0];
  _RAND_305 = {1{`RANDOM}};
  signReg_20 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  multiplierReg_21 = _RAND_306[4:0];
  _RAND_307 = {1{`RANDOM}};
  signReg_21 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  multiplierReg_22 = _RAND_308[4:0];
  _RAND_309 = {1{`RANDOM}};
  signReg_22 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  multiplierReg_23 = _RAND_310[4:0];
  _RAND_311 = {1{`RANDOM}};
  signReg_23 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  multiplierReg_24 = _RAND_312[4:0];
  _RAND_313 = {1{`RANDOM}};
  signReg_24 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  multiplierReg_25 = _RAND_314[4:0];
  _RAND_315 = {1{`RANDOM}};
  signReg_25 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  multiplierReg_26 = _RAND_316[4:0];
  _RAND_317 = {1{`RANDOM}};
  signReg_26 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  multiplierReg_27 = _RAND_318[4:0];
  _RAND_319 = {1{`RANDOM}};
  signReg_27 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  multiplierReg_28 = _RAND_320[4:0];
  _RAND_321 = {1{`RANDOM}};
  signReg_28 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  multiplierReg_29 = _RAND_322[4:0];
  _RAND_323 = {1{`RANDOM}};
  signReg_29 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  multiplierReg_30 = _RAND_324[4:0];
  _RAND_325 = {1{`RANDOM}};
  signReg_30 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  multiplierReg_31 = _RAND_326[4:0];
  _RAND_327 = {1{`RANDOM}};
  signReg_31 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  multiplierReg_32 = _RAND_328[4:0];
  _RAND_329 = {1{`RANDOM}};
  signReg_32 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  multiplierReg_33 = _RAND_330[4:0];
  _RAND_331 = {1{`RANDOM}};
  signReg_33 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  multiplierReg_34 = _RAND_332[4:0];
  _RAND_333 = {1{`RANDOM}};
  signReg_34 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  multiplierReg_35 = _RAND_334[4:0];
  _RAND_335 = {1{`RANDOM}};
  signReg_35 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  multiplierReg_36 = _RAND_336[4:0];
  _RAND_337 = {1{`RANDOM}};
  signReg_36 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  multiplierReg_37 = _RAND_338[4:0];
  _RAND_339 = {1{`RANDOM}};
  signReg_37 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  multiplierReg_38 = _RAND_340[4:0];
  _RAND_341 = {1{`RANDOM}};
  signReg_38 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  multiplierReg_39 = _RAND_342[4:0];
  _RAND_343 = {1{`RANDOM}};
  signReg_39 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  multiplierReg_40 = _RAND_344[4:0];
  _RAND_345 = {1{`RANDOM}};
  signReg_40 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  multiplierReg_41 = _RAND_346[4:0];
  _RAND_347 = {1{`RANDOM}};
  signReg_41 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  multiplierReg_42 = _RAND_348[4:0];
  _RAND_349 = {1{`RANDOM}};
  signReg_42 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  multiplierReg_43 = _RAND_350[4:0];
  _RAND_351 = {1{`RANDOM}};
  signReg_43 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  multiplierReg_44 = _RAND_352[4:0];
  _RAND_353 = {1{`RANDOM}};
  signReg_44 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  multiplierReg_45 = _RAND_354[4:0];
  _RAND_355 = {1{`RANDOM}};
  signReg_45 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  multiplierReg_46 = _RAND_356[4:0];
  _RAND_357 = {1{`RANDOM}};
  signReg_46 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  multiplierReg_47 = _RAND_358[4:0];
  _RAND_359 = {1{`RANDOM}};
  signReg_47 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  multiplierReg_48 = _RAND_360[4:0];
  _RAND_361 = {1{`RANDOM}};
  signReg_48 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  multiplierReg_49 = _RAND_362[4:0];
  _RAND_363 = {1{`RANDOM}};
  signReg_49 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  multiplierReg_50 = _RAND_364[4:0];
  _RAND_365 = {1{`RANDOM}};
  signReg_50 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  multiplierReg_51 = _RAND_366[4:0];
  _RAND_367 = {1{`RANDOM}};
  signReg_51 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  multiplierReg_52 = _RAND_368[4:0];
  _RAND_369 = {1{`RANDOM}};
  signReg_52 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  multiplierReg_53 = _RAND_370[4:0];
  _RAND_371 = {1{`RANDOM}};
  signReg_53 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  multiplierReg_54 = _RAND_372[4:0];
  _RAND_373 = {1{`RANDOM}};
  signReg_54 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  multiplierReg_55 = _RAND_374[4:0];
  _RAND_375 = {1{`RANDOM}};
  signReg_55 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  multiplierReg_56 = _RAND_376[4:0];
  _RAND_377 = {1{`RANDOM}};
  signReg_56 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  multiplierReg_57 = _RAND_378[4:0];
  _RAND_379 = {1{`RANDOM}};
  signReg_57 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  multiplierReg_58 = _RAND_380[4:0];
  _RAND_381 = {1{`RANDOM}};
  signReg_58 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  multiplierReg_59 = _RAND_382[4:0];
  _RAND_383 = {1{`RANDOM}};
  signReg_59 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  multiplierReg_60 = _RAND_384[4:0];
  _RAND_385 = {1{`RANDOM}};
  signReg_60 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  multiplierReg_61 = _RAND_386[4:0];
  _RAND_387 = {1{`RANDOM}};
  signReg_61 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  multiplierReg_62 = _RAND_388[4:0];
  _RAND_389 = {1{`RANDOM}};
  signReg_62 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  multiplierReg_63 = _RAND_390[4:0];
  _RAND_391 = {1{`RANDOM}};
  signReg_63 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  dotProductRegs_1_0 = _RAND_392[4:0];
  _RAND_393 = {1{`RANDOM}};
  dotProductRegs_1_1 = _RAND_393[4:0];
  _RAND_394 = {1{`RANDOM}};
  dotProductRegs_1_2 = _RAND_394[4:0];
  _RAND_395 = {1{`RANDOM}};
  dotProductRegs_1_3 = _RAND_395[4:0];
  _RAND_396 = {1{`RANDOM}};
  dotProductRegs_1_4 = _RAND_396[4:0];
  _RAND_397 = {1{`RANDOM}};
  dotProductRegs_1_5 = _RAND_397[4:0];
  _RAND_398 = {1{`RANDOM}};
  dotProductRegs_1_6 = _RAND_398[4:0];
  _RAND_399 = {1{`RANDOM}};
  dotProductRegs_1_7 = _RAND_399[4:0];
  _RAND_400 = {1{`RANDOM}};
  dotProductRegs_1_8 = _RAND_400[4:0];
  _RAND_401 = {1{`RANDOM}};
  dotProductRegs_1_9 = _RAND_401[4:0];
  _RAND_402 = {1{`RANDOM}};
  dotProductRegs_1_10 = _RAND_402[4:0];
  _RAND_403 = {1{`RANDOM}};
  dotProductRegs_1_11 = _RAND_403[4:0];
  _RAND_404 = {1{`RANDOM}};
  dotProductRegs_1_12 = _RAND_404[4:0];
  _RAND_405 = {1{`RANDOM}};
  dotProductRegs_1_13 = _RAND_405[4:0];
  _RAND_406 = {1{`RANDOM}};
  dotProductRegs_1_14 = _RAND_406[4:0];
  _RAND_407 = {1{`RANDOM}};
  dotProductRegs_1_15 = _RAND_407[4:0];
  _RAND_408 = {1{`RANDOM}};
  dotProductRegs_1_16 = _RAND_408[4:0];
  _RAND_409 = {1{`RANDOM}};
  dotProductRegs_1_17 = _RAND_409[4:0];
  _RAND_410 = {1{`RANDOM}};
  dotProductRegs_1_18 = _RAND_410[4:0];
  _RAND_411 = {1{`RANDOM}};
  dotProductRegs_1_19 = _RAND_411[4:0];
  _RAND_412 = {1{`RANDOM}};
  dotProductRegs_1_20 = _RAND_412[4:0];
  _RAND_413 = {1{`RANDOM}};
  dotProductRegs_1_21 = _RAND_413[4:0];
  _RAND_414 = {1{`RANDOM}};
  dotProductRegs_1_22 = _RAND_414[4:0];
  _RAND_415 = {1{`RANDOM}};
  dotProductRegs_1_23 = _RAND_415[4:0];
  _RAND_416 = {1{`RANDOM}};
  dotProductRegs_1_24 = _RAND_416[4:0];
  _RAND_417 = {1{`RANDOM}};
  dotProductRegs_1_25 = _RAND_417[4:0];
  _RAND_418 = {1{`RANDOM}};
  dotProductRegs_1_26 = _RAND_418[4:0];
  _RAND_419 = {1{`RANDOM}};
  dotProductRegs_1_27 = _RAND_419[4:0];
  _RAND_420 = {1{`RANDOM}};
  dotProductRegs_1_28 = _RAND_420[4:0];
  _RAND_421 = {1{`RANDOM}};
  dotProductRegs_1_29 = _RAND_421[4:0];
  _RAND_422 = {1{`RANDOM}};
  dotProductRegs_1_30 = _RAND_422[4:0];
  _RAND_423 = {1{`RANDOM}};
  dotProductRegs_1_31 = _RAND_423[4:0];
  _RAND_424 = {1{`RANDOM}};
  dotProductRegs_1_32 = _RAND_424[4:0];
  _RAND_425 = {1{`RANDOM}};
  dotProductRegs_1_33 = _RAND_425[4:0];
  _RAND_426 = {1{`RANDOM}};
  dotProductRegs_1_34 = _RAND_426[4:0];
  _RAND_427 = {1{`RANDOM}};
  dotProductRegs_1_35 = _RAND_427[4:0];
  _RAND_428 = {1{`RANDOM}};
  dotProductRegs_1_36 = _RAND_428[4:0];
  _RAND_429 = {1{`RANDOM}};
  dotProductRegs_1_37 = _RAND_429[4:0];
  _RAND_430 = {1{`RANDOM}};
  dotProductRegs_1_38 = _RAND_430[4:0];
  _RAND_431 = {1{`RANDOM}};
  dotProductRegs_1_39 = _RAND_431[4:0];
  _RAND_432 = {1{`RANDOM}};
  dotProductRegs_1_40 = _RAND_432[4:0];
  _RAND_433 = {1{`RANDOM}};
  dotProductRegs_1_41 = _RAND_433[4:0];
  _RAND_434 = {1{`RANDOM}};
  dotProductRegs_1_42 = _RAND_434[4:0];
  _RAND_435 = {1{`RANDOM}};
  dotProductRegs_1_43 = _RAND_435[4:0];
  _RAND_436 = {1{`RANDOM}};
  dotProductRegs_1_44 = _RAND_436[4:0];
  _RAND_437 = {1{`RANDOM}};
  dotProductRegs_1_45 = _RAND_437[4:0];
  _RAND_438 = {1{`RANDOM}};
  dotProductRegs_1_46 = _RAND_438[4:0];
  _RAND_439 = {1{`RANDOM}};
  dotProductRegs_1_47 = _RAND_439[4:0];
  _RAND_440 = {1{`RANDOM}};
  dotProductRegs_1_48 = _RAND_440[4:0];
  _RAND_441 = {1{`RANDOM}};
  dotProductRegs_1_49 = _RAND_441[4:0];
  _RAND_442 = {1{`RANDOM}};
  dotProductRegs_1_50 = _RAND_442[4:0];
  _RAND_443 = {1{`RANDOM}};
  dotProductRegs_1_51 = _RAND_443[4:0];
  _RAND_444 = {1{`RANDOM}};
  dotProductRegs_1_52 = _RAND_444[4:0];
  _RAND_445 = {1{`RANDOM}};
  dotProductRegs_1_53 = _RAND_445[4:0];
  _RAND_446 = {1{`RANDOM}};
  dotProductRegs_1_54 = _RAND_446[4:0];
  _RAND_447 = {1{`RANDOM}};
  dotProductRegs_1_55 = _RAND_447[4:0];
  _RAND_448 = {1{`RANDOM}};
  dotProductRegs_1_56 = _RAND_448[4:0];
  _RAND_449 = {1{`RANDOM}};
  dotProductRegs_1_57 = _RAND_449[4:0];
  _RAND_450 = {1{`RANDOM}};
  dotProductRegs_1_58 = _RAND_450[4:0];
  _RAND_451 = {1{`RANDOM}};
  dotProductRegs_1_59 = _RAND_451[4:0];
  _RAND_452 = {1{`RANDOM}};
  dotProductRegs_1_60 = _RAND_452[4:0];
  _RAND_453 = {1{`RANDOM}};
  dotProductRegs_1_61 = _RAND_453[4:0];
  _RAND_454 = {1{`RANDOM}};
  dotProductRegs_1_62 = _RAND_454[4:0];
  _RAND_455 = {1{`RANDOM}};
  dotProductRegs_1_63 = _RAND_455[4:0];
  _RAND_456 = {1{`RANDOM}};
  signs_1_0 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  signs_1_1 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  signs_1_2 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  signs_1_3 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  signs_1_4 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  signs_1_5 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  signs_1_6 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  signs_1_7 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  signs_1_8 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  signs_1_9 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  signs_1_10 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  signs_1_11 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  signs_1_12 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  signs_1_13 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  signs_1_14 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  signs_1_15 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  signs_1_16 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  signs_1_17 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  signs_1_18 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  signs_1_19 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  signs_1_20 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  signs_1_21 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  signs_1_22 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  signs_1_23 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  signs_1_24 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  signs_1_25 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  signs_1_26 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  signs_1_27 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  signs_1_28 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  signs_1_29 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  signs_1_30 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  signs_1_31 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  signs_1_32 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  signs_1_33 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  signs_1_34 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  signs_1_35 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  signs_1_36 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  signs_1_37 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  signs_1_38 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  signs_1_39 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  signs_1_40 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  signs_1_41 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  signs_1_42 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  signs_1_43 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  signs_1_44 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  signs_1_45 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  signs_1_46 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  signs_1_47 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  signs_1_48 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  signs_1_49 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  signs_1_50 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  signs_1_51 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  signs_1_52 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  signs_1_53 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  signs_1_54 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  signs_1_55 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  signs_1_56 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  signs_1_57 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  signs_1_58 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  signs_1_59 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  signs_1_60 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  signs_1_61 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  signs_1_62 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  signs_1_63 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  two_complement_1_0 = _RAND_520[5:0];
  _RAND_521 = {1{`RANDOM}};
  two_complement_1_1 = _RAND_521[5:0];
  _RAND_522 = {1{`RANDOM}};
  two_complement_1_2 = _RAND_522[5:0];
  _RAND_523 = {1{`RANDOM}};
  two_complement_1_3 = _RAND_523[5:0];
  _RAND_524 = {1{`RANDOM}};
  two_complement_1_4 = _RAND_524[5:0];
  _RAND_525 = {1{`RANDOM}};
  two_complement_1_5 = _RAND_525[5:0];
  _RAND_526 = {1{`RANDOM}};
  two_complement_1_6 = _RAND_526[5:0];
  _RAND_527 = {1{`RANDOM}};
  two_complement_1_7 = _RAND_527[5:0];
  _RAND_528 = {1{`RANDOM}};
  two_complement_1_8 = _RAND_528[5:0];
  _RAND_529 = {1{`RANDOM}};
  two_complement_1_9 = _RAND_529[5:0];
  _RAND_530 = {1{`RANDOM}};
  two_complement_1_10 = _RAND_530[5:0];
  _RAND_531 = {1{`RANDOM}};
  two_complement_1_11 = _RAND_531[5:0];
  _RAND_532 = {1{`RANDOM}};
  two_complement_1_12 = _RAND_532[5:0];
  _RAND_533 = {1{`RANDOM}};
  two_complement_1_13 = _RAND_533[5:0];
  _RAND_534 = {1{`RANDOM}};
  two_complement_1_14 = _RAND_534[5:0];
  _RAND_535 = {1{`RANDOM}};
  two_complement_1_15 = _RAND_535[5:0];
  _RAND_536 = {1{`RANDOM}};
  two_complement_1_16 = _RAND_536[5:0];
  _RAND_537 = {1{`RANDOM}};
  two_complement_1_17 = _RAND_537[5:0];
  _RAND_538 = {1{`RANDOM}};
  two_complement_1_18 = _RAND_538[5:0];
  _RAND_539 = {1{`RANDOM}};
  two_complement_1_19 = _RAND_539[5:0];
  _RAND_540 = {1{`RANDOM}};
  two_complement_1_20 = _RAND_540[5:0];
  _RAND_541 = {1{`RANDOM}};
  two_complement_1_21 = _RAND_541[5:0];
  _RAND_542 = {1{`RANDOM}};
  two_complement_1_22 = _RAND_542[5:0];
  _RAND_543 = {1{`RANDOM}};
  two_complement_1_23 = _RAND_543[5:0];
  _RAND_544 = {1{`RANDOM}};
  two_complement_1_24 = _RAND_544[5:0];
  _RAND_545 = {1{`RANDOM}};
  two_complement_1_25 = _RAND_545[5:0];
  _RAND_546 = {1{`RANDOM}};
  two_complement_1_26 = _RAND_546[5:0];
  _RAND_547 = {1{`RANDOM}};
  two_complement_1_27 = _RAND_547[5:0];
  _RAND_548 = {1{`RANDOM}};
  two_complement_1_28 = _RAND_548[5:0];
  _RAND_549 = {1{`RANDOM}};
  two_complement_1_29 = _RAND_549[5:0];
  _RAND_550 = {1{`RANDOM}};
  two_complement_1_30 = _RAND_550[5:0];
  _RAND_551 = {1{`RANDOM}};
  two_complement_1_31 = _RAND_551[5:0];
  _RAND_552 = {1{`RANDOM}};
  two_complement_1_32 = _RAND_552[5:0];
  _RAND_553 = {1{`RANDOM}};
  two_complement_1_33 = _RAND_553[5:0];
  _RAND_554 = {1{`RANDOM}};
  two_complement_1_34 = _RAND_554[5:0];
  _RAND_555 = {1{`RANDOM}};
  two_complement_1_35 = _RAND_555[5:0];
  _RAND_556 = {1{`RANDOM}};
  two_complement_1_36 = _RAND_556[5:0];
  _RAND_557 = {1{`RANDOM}};
  two_complement_1_37 = _RAND_557[5:0];
  _RAND_558 = {1{`RANDOM}};
  two_complement_1_38 = _RAND_558[5:0];
  _RAND_559 = {1{`RANDOM}};
  two_complement_1_39 = _RAND_559[5:0];
  _RAND_560 = {1{`RANDOM}};
  two_complement_1_40 = _RAND_560[5:0];
  _RAND_561 = {1{`RANDOM}};
  two_complement_1_41 = _RAND_561[5:0];
  _RAND_562 = {1{`RANDOM}};
  two_complement_1_42 = _RAND_562[5:0];
  _RAND_563 = {1{`RANDOM}};
  two_complement_1_43 = _RAND_563[5:0];
  _RAND_564 = {1{`RANDOM}};
  two_complement_1_44 = _RAND_564[5:0];
  _RAND_565 = {1{`RANDOM}};
  two_complement_1_45 = _RAND_565[5:0];
  _RAND_566 = {1{`RANDOM}};
  two_complement_1_46 = _RAND_566[5:0];
  _RAND_567 = {1{`RANDOM}};
  two_complement_1_47 = _RAND_567[5:0];
  _RAND_568 = {1{`RANDOM}};
  two_complement_1_48 = _RAND_568[5:0];
  _RAND_569 = {1{`RANDOM}};
  two_complement_1_49 = _RAND_569[5:0];
  _RAND_570 = {1{`RANDOM}};
  two_complement_1_50 = _RAND_570[5:0];
  _RAND_571 = {1{`RANDOM}};
  two_complement_1_51 = _RAND_571[5:0];
  _RAND_572 = {1{`RANDOM}};
  two_complement_1_52 = _RAND_572[5:0];
  _RAND_573 = {1{`RANDOM}};
  two_complement_1_53 = _RAND_573[5:0];
  _RAND_574 = {1{`RANDOM}};
  two_complement_1_54 = _RAND_574[5:0];
  _RAND_575 = {1{`RANDOM}};
  two_complement_1_55 = _RAND_575[5:0];
  _RAND_576 = {1{`RANDOM}};
  two_complement_1_56 = _RAND_576[5:0];
  _RAND_577 = {1{`RANDOM}};
  two_complement_1_57 = _RAND_577[5:0];
  _RAND_578 = {1{`RANDOM}};
  two_complement_1_58 = _RAND_578[5:0];
  _RAND_579 = {1{`RANDOM}};
  two_complement_1_59 = _RAND_579[5:0];
  _RAND_580 = {1{`RANDOM}};
  two_complement_1_60 = _RAND_580[5:0];
  _RAND_581 = {1{`RANDOM}};
  two_complement_1_61 = _RAND_581[5:0];
  _RAND_582 = {1{`RANDOM}};
  two_complement_1_62 = _RAND_582[5:0];
  _RAND_583 = {1{`RANDOM}};
  two_complement_1_63 = _RAND_583[5:0];
  _RAND_584 = {1{`RANDOM}};
  two_complement_buffer_1_0 = _RAND_584[5:0];
  _RAND_585 = {1{`RANDOM}};
  two_complement_buffer_1_1 = _RAND_585[5:0];
  _RAND_586 = {1{`RANDOM}};
  two_complement_buffer_1_2 = _RAND_586[5:0];
  _RAND_587 = {1{`RANDOM}};
  two_complement_buffer_1_3 = _RAND_587[5:0];
  _RAND_588 = {1{`RANDOM}};
  two_complement_buffer_1_4 = _RAND_588[5:0];
  _RAND_589 = {1{`RANDOM}};
  two_complement_buffer_1_5 = _RAND_589[5:0];
  _RAND_590 = {1{`RANDOM}};
  two_complement_buffer_1_6 = _RAND_590[5:0];
  _RAND_591 = {1{`RANDOM}};
  two_complement_buffer_1_7 = _RAND_591[5:0];
  _RAND_592 = {1{`RANDOM}};
  two_complement_buffer_1_8 = _RAND_592[5:0];
  _RAND_593 = {1{`RANDOM}};
  two_complement_buffer_1_9 = _RAND_593[5:0];
  _RAND_594 = {1{`RANDOM}};
  two_complement_buffer_1_10 = _RAND_594[5:0];
  _RAND_595 = {1{`RANDOM}};
  two_complement_buffer_1_11 = _RAND_595[5:0];
  _RAND_596 = {1{`RANDOM}};
  two_complement_buffer_1_12 = _RAND_596[5:0];
  _RAND_597 = {1{`RANDOM}};
  two_complement_buffer_1_13 = _RAND_597[5:0];
  _RAND_598 = {1{`RANDOM}};
  two_complement_buffer_1_14 = _RAND_598[5:0];
  _RAND_599 = {1{`RANDOM}};
  two_complement_buffer_1_15 = _RAND_599[5:0];
  _RAND_600 = {1{`RANDOM}};
  two_complement_buffer_1_16 = _RAND_600[5:0];
  _RAND_601 = {1{`RANDOM}};
  two_complement_buffer_1_17 = _RAND_601[5:0];
  _RAND_602 = {1{`RANDOM}};
  two_complement_buffer_1_18 = _RAND_602[5:0];
  _RAND_603 = {1{`RANDOM}};
  two_complement_buffer_1_19 = _RAND_603[5:0];
  _RAND_604 = {1{`RANDOM}};
  two_complement_buffer_1_20 = _RAND_604[5:0];
  _RAND_605 = {1{`RANDOM}};
  two_complement_buffer_1_21 = _RAND_605[5:0];
  _RAND_606 = {1{`RANDOM}};
  two_complement_buffer_1_22 = _RAND_606[5:0];
  _RAND_607 = {1{`RANDOM}};
  two_complement_buffer_1_23 = _RAND_607[5:0];
  _RAND_608 = {1{`RANDOM}};
  two_complement_buffer_1_24 = _RAND_608[5:0];
  _RAND_609 = {1{`RANDOM}};
  two_complement_buffer_1_25 = _RAND_609[5:0];
  _RAND_610 = {1{`RANDOM}};
  two_complement_buffer_1_26 = _RAND_610[5:0];
  _RAND_611 = {1{`RANDOM}};
  two_complement_buffer_1_27 = _RAND_611[5:0];
  _RAND_612 = {1{`RANDOM}};
  two_complement_buffer_1_28 = _RAND_612[5:0];
  _RAND_613 = {1{`RANDOM}};
  two_complement_buffer_1_29 = _RAND_613[5:0];
  _RAND_614 = {1{`RANDOM}};
  two_complement_buffer_1_30 = _RAND_614[5:0];
  _RAND_615 = {1{`RANDOM}};
  two_complement_buffer_1_31 = _RAND_615[5:0];
  _RAND_616 = {1{`RANDOM}};
  two_complement_buffer_1_32 = _RAND_616[5:0];
  _RAND_617 = {1{`RANDOM}};
  two_complement_buffer_1_33 = _RAND_617[5:0];
  _RAND_618 = {1{`RANDOM}};
  two_complement_buffer_1_34 = _RAND_618[5:0];
  _RAND_619 = {1{`RANDOM}};
  two_complement_buffer_1_35 = _RAND_619[5:0];
  _RAND_620 = {1{`RANDOM}};
  two_complement_buffer_1_36 = _RAND_620[5:0];
  _RAND_621 = {1{`RANDOM}};
  two_complement_buffer_1_37 = _RAND_621[5:0];
  _RAND_622 = {1{`RANDOM}};
  two_complement_buffer_1_38 = _RAND_622[5:0];
  _RAND_623 = {1{`RANDOM}};
  two_complement_buffer_1_39 = _RAND_623[5:0];
  _RAND_624 = {1{`RANDOM}};
  two_complement_buffer_1_40 = _RAND_624[5:0];
  _RAND_625 = {1{`RANDOM}};
  two_complement_buffer_1_41 = _RAND_625[5:0];
  _RAND_626 = {1{`RANDOM}};
  two_complement_buffer_1_42 = _RAND_626[5:0];
  _RAND_627 = {1{`RANDOM}};
  two_complement_buffer_1_43 = _RAND_627[5:0];
  _RAND_628 = {1{`RANDOM}};
  two_complement_buffer_1_44 = _RAND_628[5:0];
  _RAND_629 = {1{`RANDOM}};
  two_complement_buffer_1_45 = _RAND_629[5:0];
  _RAND_630 = {1{`RANDOM}};
  two_complement_buffer_1_46 = _RAND_630[5:0];
  _RAND_631 = {1{`RANDOM}};
  two_complement_buffer_1_47 = _RAND_631[5:0];
  _RAND_632 = {1{`RANDOM}};
  two_complement_buffer_1_48 = _RAND_632[5:0];
  _RAND_633 = {1{`RANDOM}};
  two_complement_buffer_1_49 = _RAND_633[5:0];
  _RAND_634 = {1{`RANDOM}};
  two_complement_buffer_1_50 = _RAND_634[5:0];
  _RAND_635 = {1{`RANDOM}};
  two_complement_buffer_1_51 = _RAND_635[5:0];
  _RAND_636 = {1{`RANDOM}};
  two_complement_buffer_1_52 = _RAND_636[5:0];
  _RAND_637 = {1{`RANDOM}};
  two_complement_buffer_1_53 = _RAND_637[5:0];
  _RAND_638 = {1{`RANDOM}};
  two_complement_buffer_1_54 = _RAND_638[5:0];
  _RAND_639 = {1{`RANDOM}};
  two_complement_buffer_1_55 = _RAND_639[5:0];
  _RAND_640 = {1{`RANDOM}};
  two_complement_buffer_1_56 = _RAND_640[5:0];
  _RAND_641 = {1{`RANDOM}};
  two_complement_buffer_1_57 = _RAND_641[5:0];
  _RAND_642 = {1{`RANDOM}};
  two_complement_buffer_1_58 = _RAND_642[5:0];
  _RAND_643 = {1{`RANDOM}};
  two_complement_buffer_1_59 = _RAND_643[5:0];
  _RAND_644 = {1{`RANDOM}};
  two_complement_buffer_1_60 = _RAND_644[5:0];
  _RAND_645 = {1{`RANDOM}};
  two_complement_buffer_1_61 = _RAND_645[5:0];
  _RAND_646 = {1{`RANDOM}};
  two_complement_buffer_1_62 = _RAND_646[5:0];
  _RAND_647 = {1{`RANDOM}};
  two_complement_buffer_1_63 = _RAND_647[5:0];
  _RAND_648 = {1{`RANDOM}};
  multiplierReg_64 = _RAND_648[4:0];
  _RAND_649 = {1{`RANDOM}};
  signReg_64 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  multiplierReg_65 = _RAND_650[4:0];
  _RAND_651 = {1{`RANDOM}};
  signReg_65 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  multiplierReg_66 = _RAND_652[4:0];
  _RAND_653 = {1{`RANDOM}};
  signReg_66 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  multiplierReg_67 = _RAND_654[4:0];
  _RAND_655 = {1{`RANDOM}};
  signReg_67 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  multiplierReg_68 = _RAND_656[4:0];
  _RAND_657 = {1{`RANDOM}};
  signReg_68 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  multiplierReg_69 = _RAND_658[4:0];
  _RAND_659 = {1{`RANDOM}};
  signReg_69 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  multiplierReg_70 = _RAND_660[4:0];
  _RAND_661 = {1{`RANDOM}};
  signReg_70 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  multiplierReg_71 = _RAND_662[4:0];
  _RAND_663 = {1{`RANDOM}};
  signReg_71 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  multiplierReg_72 = _RAND_664[4:0];
  _RAND_665 = {1{`RANDOM}};
  signReg_72 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  multiplierReg_73 = _RAND_666[4:0];
  _RAND_667 = {1{`RANDOM}};
  signReg_73 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  multiplierReg_74 = _RAND_668[4:0];
  _RAND_669 = {1{`RANDOM}};
  signReg_74 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  multiplierReg_75 = _RAND_670[4:0];
  _RAND_671 = {1{`RANDOM}};
  signReg_75 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  multiplierReg_76 = _RAND_672[4:0];
  _RAND_673 = {1{`RANDOM}};
  signReg_76 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  multiplierReg_77 = _RAND_674[4:0];
  _RAND_675 = {1{`RANDOM}};
  signReg_77 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  multiplierReg_78 = _RAND_676[4:0];
  _RAND_677 = {1{`RANDOM}};
  signReg_78 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  multiplierReg_79 = _RAND_678[4:0];
  _RAND_679 = {1{`RANDOM}};
  signReg_79 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  multiplierReg_80 = _RAND_680[4:0];
  _RAND_681 = {1{`RANDOM}};
  signReg_80 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  multiplierReg_81 = _RAND_682[4:0];
  _RAND_683 = {1{`RANDOM}};
  signReg_81 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  multiplierReg_82 = _RAND_684[4:0];
  _RAND_685 = {1{`RANDOM}};
  signReg_82 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  multiplierReg_83 = _RAND_686[4:0];
  _RAND_687 = {1{`RANDOM}};
  signReg_83 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  multiplierReg_84 = _RAND_688[4:0];
  _RAND_689 = {1{`RANDOM}};
  signReg_84 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  multiplierReg_85 = _RAND_690[4:0];
  _RAND_691 = {1{`RANDOM}};
  signReg_85 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  multiplierReg_86 = _RAND_692[4:0];
  _RAND_693 = {1{`RANDOM}};
  signReg_86 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  multiplierReg_87 = _RAND_694[4:0];
  _RAND_695 = {1{`RANDOM}};
  signReg_87 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  multiplierReg_88 = _RAND_696[4:0];
  _RAND_697 = {1{`RANDOM}};
  signReg_88 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  multiplierReg_89 = _RAND_698[4:0];
  _RAND_699 = {1{`RANDOM}};
  signReg_89 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  multiplierReg_90 = _RAND_700[4:0];
  _RAND_701 = {1{`RANDOM}};
  signReg_90 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  multiplierReg_91 = _RAND_702[4:0];
  _RAND_703 = {1{`RANDOM}};
  signReg_91 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  multiplierReg_92 = _RAND_704[4:0];
  _RAND_705 = {1{`RANDOM}};
  signReg_92 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  multiplierReg_93 = _RAND_706[4:0];
  _RAND_707 = {1{`RANDOM}};
  signReg_93 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  multiplierReg_94 = _RAND_708[4:0];
  _RAND_709 = {1{`RANDOM}};
  signReg_94 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  multiplierReg_95 = _RAND_710[4:0];
  _RAND_711 = {1{`RANDOM}};
  signReg_95 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  multiplierReg_96 = _RAND_712[4:0];
  _RAND_713 = {1{`RANDOM}};
  signReg_96 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  multiplierReg_97 = _RAND_714[4:0];
  _RAND_715 = {1{`RANDOM}};
  signReg_97 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  multiplierReg_98 = _RAND_716[4:0];
  _RAND_717 = {1{`RANDOM}};
  signReg_98 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  multiplierReg_99 = _RAND_718[4:0];
  _RAND_719 = {1{`RANDOM}};
  signReg_99 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  multiplierReg_100 = _RAND_720[4:0];
  _RAND_721 = {1{`RANDOM}};
  signReg_100 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  multiplierReg_101 = _RAND_722[4:0];
  _RAND_723 = {1{`RANDOM}};
  signReg_101 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  multiplierReg_102 = _RAND_724[4:0];
  _RAND_725 = {1{`RANDOM}};
  signReg_102 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  multiplierReg_103 = _RAND_726[4:0];
  _RAND_727 = {1{`RANDOM}};
  signReg_103 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  multiplierReg_104 = _RAND_728[4:0];
  _RAND_729 = {1{`RANDOM}};
  signReg_104 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  multiplierReg_105 = _RAND_730[4:0];
  _RAND_731 = {1{`RANDOM}};
  signReg_105 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  multiplierReg_106 = _RAND_732[4:0];
  _RAND_733 = {1{`RANDOM}};
  signReg_106 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  multiplierReg_107 = _RAND_734[4:0];
  _RAND_735 = {1{`RANDOM}};
  signReg_107 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  multiplierReg_108 = _RAND_736[4:0];
  _RAND_737 = {1{`RANDOM}};
  signReg_108 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  multiplierReg_109 = _RAND_738[4:0];
  _RAND_739 = {1{`RANDOM}};
  signReg_109 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  multiplierReg_110 = _RAND_740[4:0];
  _RAND_741 = {1{`RANDOM}};
  signReg_110 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  multiplierReg_111 = _RAND_742[4:0];
  _RAND_743 = {1{`RANDOM}};
  signReg_111 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  multiplierReg_112 = _RAND_744[4:0];
  _RAND_745 = {1{`RANDOM}};
  signReg_112 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  multiplierReg_113 = _RAND_746[4:0];
  _RAND_747 = {1{`RANDOM}};
  signReg_113 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  multiplierReg_114 = _RAND_748[4:0];
  _RAND_749 = {1{`RANDOM}};
  signReg_114 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  multiplierReg_115 = _RAND_750[4:0];
  _RAND_751 = {1{`RANDOM}};
  signReg_115 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  multiplierReg_116 = _RAND_752[4:0];
  _RAND_753 = {1{`RANDOM}};
  signReg_116 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  multiplierReg_117 = _RAND_754[4:0];
  _RAND_755 = {1{`RANDOM}};
  signReg_117 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  multiplierReg_118 = _RAND_756[4:0];
  _RAND_757 = {1{`RANDOM}};
  signReg_118 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  multiplierReg_119 = _RAND_758[4:0];
  _RAND_759 = {1{`RANDOM}};
  signReg_119 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  multiplierReg_120 = _RAND_760[4:0];
  _RAND_761 = {1{`RANDOM}};
  signReg_120 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  multiplierReg_121 = _RAND_762[4:0];
  _RAND_763 = {1{`RANDOM}};
  signReg_121 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  multiplierReg_122 = _RAND_764[4:0];
  _RAND_765 = {1{`RANDOM}};
  signReg_122 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  multiplierReg_123 = _RAND_766[4:0];
  _RAND_767 = {1{`RANDOM}};
  signReg_123 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  multiplierReg_124 = _RAND_768[4:0];
  _RAND_769 = {1{`RANDOM}};
  signReg_124 = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  multiplierReg_125 = _RAND_770[4:0];
  _RAND_771 = {1{`RANDOM}};
  signReg_125 = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  multiplierReg_126 = _RAND_772[4:0];
  _RAND_773 = {1{`RANDOM}};
  signReg_126 = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  multiplierReg_127 = _RAND_774[4:0];
  _RAND_775 = {1{`RANDOM}};
  signReg_127 = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  dotProductRegs_2_0 = _RAND_776[4:0];
  _RAND_777 = {1{`RANDOM}};
  dotProductRegs_2_1 = _RAND_777[4:0];
  _RAND_778 = {1{`RANDOM}};
  dotProductRegs_2_2 = _RAND_778[4:0];
  _RAND_779 = {1{`RANDOM}};
  dotProductRegs_2_3 = _RAND_779[4:0];
  _RAND_780 = {1{`RANDOM}};
  dotProductRegs_2_4 = _RAND_780[4:0];
  _RAND_781 = {1{`RANDOM}};
  dotProductRegs_2_5 = _RAND_781[4:0];
  _RAND_782 = {1{`RANDOM}};
  dotProductRegs_2_6 = _RAND_782[4:0];
  _RAND_783 = {1{`RANDOM}};
  dotProductRegs_2_7 = _RAND_783[4:0];
  _RAND_784 = {1{`RANDOM}};
  dotProductRegs_2_8 = _RAND_784[4:0];
  _RAND_785 = {1{`RANDOM}};
  dotProductRegs_2_9 = _RAND_785[4:0];
  _RAND_786 = {1{`RANDOM}};
  dotProductRegs_2_10 = _RAND_786[4:0];
  _RAND_787 = {1{`RANDOM}};
  dotProductRegs_2_11 = _RAND_787[4:0];
  _RAND_788 = {1{`RANDOM}};
  dotProductRegs_2_12 = _RAND_788[4:0];
  _RAND_789 = {1{`RANDOM}};
  dotProductRegs_2_13 = _RAND_789[4:0];
  _RAND_790 = {1{`RANDOM}};
  dotProductRegs_2_14 = _RAND_790[4:0];
  _RAND_791 = {1{`RANDOM}};
  dotProductRegs_2_15 = _RAND_791[4:0];
  _RAND_792 = {1{`RANDOM}};
  dotProductRegs_2_16 = _RAND_792[4:0];
  _RAND_793 = {1{`RANDOM}};
  dotProductRegs_2_17 = _RAND_793[4:0];
  _RAND_794 = {1{`RANDOM}};
  dotProductRegs_2_18 = _RAND_794[4:0];
  _RAND_795 = {1{`RANDOM}};
  dotProductRegs_2_19 = _RAND_795[4:0];
  _RAND_796 = {1{`RANDOM}};
  dotProductRegs_2_20 = _RAND_796[4:0];
  _RAND_797 = {1{`RANDOM}};
  dotProductRegs_2_21 = _RAND_797[4:0];
  _RAND_798 = {1{`RANDOM}};
  dotProductRegs_2_22 = _RAND_798[4:0];
  _RAND_799 = {1{`RANDOM}};
  dotProductRegs_2_23 = _RAND_799[4:0];
  _RAND_800 = {1{`RANDOM}};
  dotProductRegs_2_24 = _RAND_800[4:0];
  _RAND_801 = {1{`RANDOM}};
  dotProductRegs_2_25 = _RAND_801[4:0];
  _RAND_802 = {1{`RANDOM}};
  dotProductRegs_2_26 = _RAND_802[4:0];
  _RAND_803 = {1{`RANDOM}};
  dotProductRegs_2_27 = _RAND_803[4:0];
  _RAND_804 = {1{`RANDOM}};
  dotProductRegs_2_28 = _RAND_804[4:0];
  _RAND_805 = {1{`RANDOM}};
  dotProductRegs_2_29 = _RAND_805[4:0];
  _RAND_806 = {1{`RANDOM}};
  dotProductRegs_2_30 = _RAND_806[4:0];
  _RAND_807 = {1{`RANDOM}};
  dotProductRegs_2_31 = _RAND_807[4:0];
  _RAND_808 = {1{`RANDOM}};
  dotProductRegs_2_32 = _RAND_808[4:0];
  _RAND_809 = {1{`RANDOM}};
  dotProductRegs_2_33 = _RAND_809[4:0];
  _RAND_810 = {1{`RANDOM}};
  dotProductRegs_2_34 = _RAND_810[4:0];
  _RAND_811 = {1{`RANDOM}};
  dotProductRegs_2_35 = _RAND_811[4:0];
  _RAND_812 = {1{`RANDOM}};
  dotProductRegs_2_36 = _RAND_812[4:0];
  _RAND_813 = {1{`RANDOM}};
  dotProductRegs_2_37 = _RAND_813[4:0];
  _RAND_814 = {1{`RANDOM}};
  dotProductRegs_2_38 = _RAND_814[4:0];
  _RAND_815 = {1{`RANDOM}};
  dotProductRegs_2_39 = _RAND_815[4:0];
  _RAND_816 = {1{`RANDOM}};
  dotProductRegs_2_40 = _RAND_816[4:0];
  _RAND_817 = {1{`RANDOM}};
  dotProductRegs_2_41 = _RAND_817[4:0];
  _RAND_818 = {1{`RANDOM}};
  dotProductRegs_2_42 = _RAND_818[4:0];
  _RAND_819 = {1{`RANDOM}};
  dotProductRegs_2_43 = _RAND_819[4:0];
  _RAND_820 = {1{`RANDOM}};
  dotProductRegs_2_44 = _RAND_820[4:0];
  _RAND_821 = {1{`RANDOM}};
  dotProductRegs_2_45 = _RAND_821[4:0];
  _RAND_822 = {1{`RANDOM}};
  dotProductRegs_2_46 = _RAND_822[4:0];
  _RAND_823 = {1{`RANDOM}};
  dotProductRegs_2_47 = _RAND_823[4:0];
  _RAND_824 = {1{`RANDOM}};
  dotProductRegs_2_48 = _RAND_824[4:0];
  _RAND_825 = {1{`RANDOM}};
  dotProductRegs_2_49 = _RAND_825[4:0];
  _RAND_826 = {1{`RANDOM}};
  dotProductRegs_2_50 = _RAND_826[4:0];
  _RAND_827 = {1{`RANDOM}};
  dotProductRegs_2_51 = _RAND_827[4:0];
  _RAND_828 = {1{`RANDOM}};
  dotProductRegs_2_52 = _RAND_828[4:0];
  _RAND_829 = {1{`RANDOM}};
  dotProductRegs_2_53 = _RAND_829[4:0];
  _RAND_830 = {1{`RANDOM}};
  dotProductRegs_2_54 = _RAND_830[4:0];
  _RAND_831 = {1{`RANDOM}};
  dotProductRegs_2_55 = _RAND_831[4:0];
  _RAND_832 = {1{`RANDOM}};
  dotProductRegs_2_56 = _RAND_832[4:0];
  _RAND_833 = {1{`RANDOM}};
  dotProductRegs_2_57 = _RAND_833[4:0];
  _RAND_834 = {1{`RANDOM}};
  dotProductRegs_2_58 = _RAND_834[4:0];
  _RAND_835 = {1{`RANDOM}};
  dotProductRegs_2_59 = _RAND_835[4:0];
  _RAND_836 = {1{`RANDOM}};
  dotProductRegs_2_60 = _RAND_836[4:0];
  _RAND_837 = {1{`RANDOM}};
  dotProductRegs_2_61 = _RAND_837[4:0];
  _RAND_838 = {1{`RANDOM}};
  dotProductRegs_2_62 = _RAND_838[4:0];
  _RAND_839 = {1{`RANDOM}};
  dotProductRegs_2_63 = _RAND_839[4:0];
  _RAND_840 = {1{`RANDOM}};
  signs_2_0 = _RAND_840[0:0];
  _RAND_841 = {1{`RANDOM}};
  signs_2_1 = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  signs_2_2 = _RAND_842[0:0];
  _RAND_843 = {1{`RANDOM}};
  signs_2_3 = _RAND_843[0:0];
  _RAND_844 = {1{`RANDOM}};
  signs_2_4 = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  signs_2_5 = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  signs_2_6 = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  signs_2_7 = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  signs_2_8 = _RAND_848[0:0];
  _RAND_849 = {1{`RANDOM}};
  signs_2_9 = _RAND_849[0:0];
  _RAND_850 = {1{`RANDOM}};
  signs_2_10 = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  signs_2_11 = _RAND_851[0:0];
  _RAND_852 = {1{`RANDOM}};
  signs_2_12 = _RAND_852[0:0];
  _RAND_853 = {1{`RANDOM}};
  signs_2_13 = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  signs_2_14 = _RAND_854[0:0];
  _RAND_855 = {1{`RANDOM}};
  signs_2_15 = _RAND_855[0:0];
  _RAND_856 = {1{`RANDOM}};
  signs_2_16 = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  signs_2_17 = _RAND_857[0:0];
  _RAND_858 = {1{`RANDOM}};
  signs_2_18 = _RAND_858[0:0];
  _RAND_859 = {1{`RANDOM}};
  signs_2_19 = _RAND_859[0:0];
  _RAND_860 = {1{`RANDOM}};
  signs_2_20 = _RAND_860[0:0];
  _RAND_861 = {1{`RANDOM}};
  signs_2_21 = _RAND_861[0:0];
  _RAND_862 = {1{`RANDOM}};
  signs_2_22 = _RAND_862[0:0];
  _RAND_863 = {1{`RANDOM}};
  signs_2_23 = _RAND_863[0:0];
  _RAND_864 = {1{`RANDOM}};
  signs_2_24 = _RAND_864[0:0];
  _RAND_865 = {1{`RANDOM}};
  signs_2_25 = _RAND_865[0:0];
  _RAND_866 = {1{`RANDOM}};
  signs_2_26 = _RAND_866[0:0];
  _RAND_867 = {1{`RANDOM}};
  signs_2_27 = _RAND_867[0:0];
  _RAND_868 = {1{`RANDOM}};
  signs_2_28 = _RAND_868[0:0];
  _RAND_869 = {1{`RANDOM}};
  signs_2_29 = _RAND_869[0:0];
  _RAND_870 = {1{`RANDOM}};
  signs_2_30 = _RAND_870[0:0];
  _RAND_871 = {1{`RANDOM}};
  signs_2_31 = _RAND_871[0:0];
  _RAND_872 = {1{`RANDOM}};
  signs_2_32 = _RAND_872[0:0];
  _RAND_873 = {1{`RANDOM}};
  signs_2_33 = _RAND_873[0:0];
  _RAND_874 = {1{`RANDOM}};
  signs_2_34 = _RAND_874[0:0];
  _RAND_875 = {1{`RANDOM}};
  signs_2_35 = _RAND_875[0:0];
  _RAND_876 = {1{`RANDOM}};
  signs_2_36 = _RAND_876[0:0];
  _RAND_877 = {1{`RANDOM}};
  signs_2_37 = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  signs_2_38 = _RAND_878[0:0];
  _RAND_879 = {1{`RANDOM}};
  signs_2_39 = _RAND_879[0:0];
  _RAND_880 = {1{`RANDOM}};
  signs_2_40 = _RAND_880[0:0];
  _RAND_881 = {1{`RANDOM}};
  signs_2_41 = _RAND_881[0:0];
  _RAND_882 = {1{`RANDOM}};
  signs_2_42 = _RAND_882[0:0];
  _RAND_883 = {1{`RANDOM}};
  signs_2_43 = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  signs_2_44 = _RAND_884[0:0];
  _RAND_885 = {1{`RANDOM}};
  signs_2_45 = _RAND_885[0:0];
  _RAND_886 = {1{`RANDOM}};
  signs_2_46 = _RAND_886[0:0];
  _RAND_887 = {1{`RANDOM}};
  signs_2_47 = _RAND_887[0:0];
  _RAND_888 = {1{`RANDOM}};
  signs_2_48 = _RAND_888[0:0];
  _RAND_889 = {1{`RANDOM}};
  signs_2_49 = _RAND_889[0:0];
  _RAND_890 = {1{`RANDOM}};
  signs_2_50 = _RAND_890[0:0];
  _RAND_891 = {1{`RANDOM}};
  signs_2_51 = _RAND_891[0:0];
  _RAND_892 = {1{`RANDOM}};
  signs_2_52 = _RAND_892[0:0];
  _RAND_893 = {1{`RANDOM}};
  signs_2_53 = _RAND_893[0:0];
  _RAND_894 = {1{`RANDOM}};
  signs_2_54 = _RAND_894[0:0];
  _RAND_895 = {1{`RANDOM}};
  signs_2_55 = _RAND_895[0:0];
  _RAND_896 = {1{`RANDOM}};
  signs_2_56 = _RAND_896[0:0];
  _RAND_897 = {1{`RANDOM}};
  signs_2_57 = _RAND_897[0:0];
  _RAND_898 = {1{`RANDOM}};
  signs_2_58 = _RAND_898[0:0];
  _RAND_899 = {1{`RANDOM}};
  signs_2_59 = _RAND_899[0:0];
  _RAND_900 = {1{`RANDOM}};
  signs_2_60 = _RAND_900[0:0];
  _RAND_901 = {1{`RANDOM}};
  signs_2_61 = _RAND_901[0:0];
  _RAND_902 = {1{`RANDOM}};
  signs_2_62 = _RAND_902[0:0];
  _RAND_903 = {1{`RANDOM}};
  signs_2_63 = _RAND_903[0:0];
  _RAND_904 = {1{`RANDOM}};
  two_complement_2_0 = _RAND_904[5:0];
  _RAND_905 = {1{`RANDOM}};
  two_complement_2_1 = _RAND_905[5:0];
  _RAND_906 = {1{`RANDOM}};
  two_complement_2_2 = _RAND_906[5:0];
  _RAND_907 = {1{`RANDOM}};
  two_complement_2_3 = _RAND_907[5:0];
  _RAND_908 = {1{`RANDOM}};
  two_complement_2_4 = _RAND_908[5:0];
  _RAND_909 = {1{`RANDOM}};
  two_complement_2_5 = _RAND_909[5:0];
  _RAND_910 = {1{`RANDOM}};
  two_complement_2_6 = _RAND_910[5:0];
  _RAND_911 = {1{`RANDOM}};
  two_complement_2_7 = _RAND_911[5:0];
  _RAND_912 = {1{`RANDOM}};
  two_complement_2_8 = _RAND_912[5:0];
  _RAND_913 = {1{`RANDOM}};
  two_complement_2_9 = _RAND_913[5:0];
  _RAND_914 = {1{`RANDOM}};
  two_complement_2_10 = _RAND_914[5:0];
  _RAND_915 = {1{`RANDOM}};
  two_complement_2_11 = _RAND_915[5:0];
  _RAND_916 = {1{`RANDOM}};
  two_complement_2_12 = _RAND_916[5:0];
  _RAND_917 = {1{`RANDOM}};
  two_complement_2_13 = _RAND_917[5:0];
  _RAND_918 = {1{`RANDOM}};
  two_complement_2_14 = _RAND_918[5:0];
  _RAND_919 = {1{`RANDOM}};
  two_complement_2_15 = _RAND_919[5:0];
  _RAND_920 = {1{`RANDOM}};
  two_complement_2_16 = _RAND_920[5:0];
  _RAND_921 = {1{`RANDOM}};
  two_complement_2_17 = _RAND_921[5:0];
  _RAND_922 = {1{`RANDOM}};
  two_complement_2_18 = _RAND_922[5:0];
  _RAND_923 = {1{`RANDOM}};
  two_complement_2_19 = _RAND_923[5:0];
  _RAND_924 = {1{`RANDOM}};
  two_complement_2_20 = _RAND_924[5:0];
  _RAND_925 = {1{`RANDOM}};
  two_complement_2_21 = _RAND_925[5:0];
  _RAND_926 = {1{`RANDOM}};
  two_complement_2_22 = _RAND_926[5:0];
  _RAND_927 = {1{`RANDOM}};
  two_complement_2_23 = _RAND_927[5:0];
  _RAND_928 = {1{`RANDOM}};
  two_complement_2_24 = _RAND_928[5:0];
  _RAND_929 = {1{`RANDOM}};
  two_complement_2_25 = _RAND_929[5:0];
  _RAND_930 = {1{`RANDOM}};
  two_complement_2_26 = _RAND_930[5:0];
  _RAND_931 = {1{`RANDOM}};
  two_complement_2_27 = _RAND_931[5:0];
  _RAND_932 = {1{`RANDOM}};
  two_complement_2_28 = _RAND_932[5:0];
  _RAND_933 = {1{`RANDOM}};
  two_complement_2_29 = _RAND_933[5:0];
  _RAND_934 = {1{`RANDOM}};
  two_complement_2_30 = _RAND_934[5:0];
  _RAND_935 = {1{`RANDOM}};
  two_complement_2_31 = _RAND_935[5:0];
  _RAND_936 = {1{`RANDOM}};
  two_complement_2_32 = _RAND_936[5:0];
  _RAND_937 = {1{`RANDOM}};
  two_complement_2_33 = _RAND_937[5:0];
  _RAND_938 = {1{`RANDOM}};
  two_complement_2_34 = _RAND_938[5:0];
  _RAND_939 = {1{`RANDOM}};
  two_complement_2_35 = _RAND_939[5:0];
  _RAND_940 = {1{`RANDOM}};
  two_complement_2_36 = _RAND_940[5:0];
  _RAND_941 = {1{`RANDOM}};
  two_complement_2_37 = _RAND_941[5:0];
  _RAND_942 = {1{`RANDOM}};
  two_complement_2_38 = _RAND_942[5:0];
  _RAND_943 = {1{`RANDOM}};
  two_complement_2_39 = _RAND_943[5:0];
  _RAND_944 = {1{`RANDOM}};
  two_complement_2_40 = _RAND_944[5:0];
  _RAND_945 = {1{`RANDOM}};
  two_complement_2_41 = _RAND_945[5:0];
  _RAND_946 = {1{`RANDOM}};
  two_complement_2_42 = _RAND_946[5:0];
  _RAND_947 = {1{`RANDOM}};
  two_complement_2_43 = _RAND_947[5:0];
  _RAND_948 = {1{`RANDOM}};
  two_complement_2_44 = _RAND_948[5:0];
  _RAND_949 = {1{`RANDOM}};
  two_complement_2_45 = _RAND_949[5:0];
  _RAND_950 = {1{`RANDOM}};
  two_complement_2_46 = _RAND_950[5:0];
  _RAND_951 = {1{`RANDOM}};
  two_complement_2_47 = _RAND_951[5:0];
  _RAND_952 = {1{`RANDOM}};
  two_complement_2_48 = _RAND_952[5:0];
  _RAND_953 = {1{`RANDOM}};
  two_complement_2_49 = _RAND_953[5:0];
  _RAND_954 = {1{`RANDOM}};
  two_complement_2_50 = _RAND_954[5:0];
  _RAND_955 = {1{`RANDOM}};
  two_complement_2_51 = _RAND_955[5:0];
  _RAND_956 = {1{`RANDOM}};
  two_complement_2_52 = _RAND_956[5:0];
  _RAND_957 = {1{`RANDOM}};
  two_complement_2_53 = _RAND_957[5:0];
  _RAND_958 = {1{`RANDOM}};
  two_complement_2_54 = _RAND_958[5:0];
  _RAND_959 = {1{`RANDOM}};
  two_complement_2_55 = _RAND_959[5:0];
  _RAND_960 = {1{`RANDOM}};
  two_complement_2_56 = _RAND_960[5:0];
  _RAND_961 = {1{`RANDOM}};
  two_complement_2_57 = _RAND_961[5:0];
  _RAND_962 = {1{`RANDOM}};
  two_complement_2_58 = _RAND_962[5:0];
  _RAND_963 = {1{`RANDOM}};
  two_complement_2_59 = _RAND_963[5:0];
  _RAND_964 = {1{`RANDOM}};
  two_complement_2_60 = _RAND_964[5:0];
  _RAND_965 = {1{`RANDOM}};
  two_complement_2_61 = _RAND_965[5:0];
  _RAND_966 = {1{`RANDOM}};
  two_complement_2_62 = _RAND_966[5:0];
  _RAND_967 = {1{`RANDOM}};
  two_complement_2_63 = _RAND_967[5:0];
  _RAND_968 = {1{`RANDOM}};
  two_complement_buffer_2_0 = _RAND_968[5:0];
  _RAND_969 = {1{`RANDOM}};
  two_complement_buffer_2_1 = _RAND_969[5:0];
  _RAND_970 = {1{`RANDOM}};
  two_complement_buffer_2_2 = _RAND_970[5:0];
  _RAND_971 = {1{`RANDOM}};
  two_complement_buffer_2_3 = _RAND_971[5:0];
  _RAND_972 = {1{`RANDOM}};
  two_complement_buffer_2_4 = _RAND_972[5:0];
  _RAND_973 = {1{`RANDOM}};
  two_complement_buffer_2_5 = _RAND_973[5:0];
  _RAND_974 = {1{`RANDOM}};
  two_complement_buffer_2_6 = _RAND_974[5:0];
  _RAND_975 = {1{`RANDOM}};
  two_complement_buffer_2_7 = _RAND_975[5:0];
  _RAND_976 = {1{`RANDOM}};
  two_complement_buffer_2_8 = _RAND_976[5:0];
  _RAND_977 = {1{`RANDOM}};
  two_complement_buffer_2_9 = _RAND_977[5:0];
  _RAND_978 = {1{`RANDOM}};
  two_complement_buffer_2_10 = _RAND_978[5:0];
  _RAND_979 = {1{`RANDOM}};
  two_complement_buffer_2_11 = _RAND_979[5:0];
  _RAND_980 = {1{`RANDOM}};
  two_complement_buffer_2_12 = _RAND_980[5:0];
  _RAND_981 = {1{`RANDOM}};
  two_complement_buffer_2_13 = _RAND_981[5:0];
  _RAND_982 = {1{`RANDOM}};
  two_complement_buffer_2_14 = _RAND_982[5:0];
  _RAND_983 = {1{`RANDOM}};
  two_complement_buffer_2_15 = _RAND_983[5:0];
  _RAND_984 = {1{`RANDOM}};
  two_complement_buffer_2_16 = _RAND_984[5:0];
  _RAND_985 = {1{`RANDOM}};
  two_complement_buffer_2_17 = _RAND_985[5:0];
  _RAND_986 = {1{`RANDOM}};
  two_complement_buffer_2_18 = _RAND_986[5:0];
  _RAND_987 = {1{`RANDOM}};
  two_complement_buffer_2_19 = _RAND_987[5:0];
  _RAND_988 = {1{`RANDOM}};
  two_complement_buffer_2_20 = _RAND_988[5:0];
  _RAND_989 = {1{`RANDOM}};
  two_complement_buffer_2_21 = _RAND_989[5:0];
  _RAND_990 = {1{`RANDOM}};
  two_complement_buffer_2_22 = _RAND_990[5:0];
  _RAND_991 = {1{`RANDOM}};
  two_complement_buffer_2_23 = _RAND_991[5:0];
  _RAND_992 = {1{`RANDOM}};
  two_complement_buffer_2_24 = _RAND_992[5:0];
  _RAND_993 = {1{`RANDOM}};
  two_complement_buffer_2_25 = _RAND_993[5:0];
  _RAND_994 = {1{`RANDOM}};
  two_complement_buffer_2_26 = _RAND_994[5:0];
  _RAND_995 = {1{`RANDOM}};
  two_complement_buffer_2_27 = _RAND_995[5:0];
  _RAND_996 = {1{`RANDOM}};
  two_complement_buffer_2_28 = _RAND_996[5:0];
  _RAND_997 = {1{`RANDOM}};
  two_complement_buffer_2_29 = _RAND_997[5:0];
  _RAND_998 = {1{`RANDOM}};
  two_complement_buffer_2_30 = _RAND_998[5:0];
  _RAND_999 = {1{`RANDOM}};
  two_complement_buffer_2_31 = _RAND_999[5:0];
  _RAND_1000 = {1{`RANDOM}};
  two_complement_buffer_2_32 = _RAND_1000[5:0];
  _RAND_1001 = {1{`RANDOM}};
  two_complement_buffer_2_33 = _RAND_1001[5:0];
  _RAND_1002 = {1{`RANDOM}};
  two_complement_buffer_2_34 = _RAND_1002[5:0];
  _RAND_1003 = {1{`RANDOM}};
  two_complement_buffer_2_35 = _RAND_1003[5:0];
  _RAND_1004 = {1{`RANDOM}};
  two_complement_buffer_2_36 = _RAND_1004[5:0];
  _RAND_1005 = {1{`RANDOM}};
  two_complement_buffer_2_37 = _RAND_1005[5:0];
  _RAND_1006 = {1{`RANDOM}};
  two_complement_buffer_2_38 = _RAND_1006[5:0];
  _RAND_1007 = {1{`RANDOM}};
  two_complement_buffer_2_39 = _RAND_1007[5:0];
  _RAND_1008 = {1{`RANDOM}};
  two_complement_buffer_2_40 = _RAND_1008[5:0];
  _RAND_1009 = {1{`RANDOM}};
  two_complement_buffer_2_41 = _RAND_1009[5:0];
  _RAND_1010 = {1{`RANDOM}};
  two_complement_buffer_2_42 = _RAND_1010[5:0];
  _RAND_1011 = {1{`RANDOM}};
  two_complement_buffer_2_43 = _RAND_1011[5:0];
  _RAND_1012 = {1{`RANDOM}};
  two_complement_buffer_2_44 = _RAND_1012[5:0];
  _RAND_1013 = {1{`RANDOM}};
  two_complement_buffer_2_45 = _RAND_1013[5:0];
  _RAND_1014 = {1{`RANDOM}};
  two_complement_buffer_2_46 = _RAND_1014[5:0];
  _RAND_1015 = {1{`RANDOM}};
  two_complement_buffer_2_47 = _RAND_1015[5:0];
  _RAND_1016 = {1{`RANDOM}};
  two_complement_buffer_2_48 = _RAND_1016[5:0];
  _RAND_1017 = {1{`RANDOM}};
  two_complement_buffer_2_49 = _RAND_1017[5:0];
  _RAND_1018 = {1{`RANDOM}};
  two_complement_buffer_2_50 = _RAND_1018[5:0];
  _RAND_1019 = {1{`RANDOM}};
  two_complement_buffer_2_51 = _RAND_1019[5:0];
  _RAND_1020 = {1{`RANDOM}};
  two_complement_buffer_2_52 = _RAND_1020[5:0];
  _RAND_1021 = {1{`RANDOM}};
  two_complement_buffer_2_53 = _RAND_1021[5:0];
  _RAND_1022 = {1{`RANDOM}};
  two_complement_buffer_2_54 = _RAND_1022[5:0];
  _RAND_1023 = {1{`RANDOM}};
  two_complement_buffer_2_55 = _RAND_1023[5:0];
  _RAND_1024 = {1{`RANDOM}};
  two_complement_buffer_2_56 = _RAND_1024[5:0];
  _RAND_1025 = {1{`RANDOM}};
  two_complement_buffer_2_57 = _RAND_1025[5:0];
  _RAND_1026 = {1{`RANDOM}};
  two_complement_buffer_2_58 = _RAND_1026[5:0];
  _RAND_1027 = {1{`RANDOM}};
  two_complement_buffer_2_59 = _RAND_1027[5:0];
  _RAND_1028 = {1{`RANDOM}};
  two_complement_buffer_2_60 = _RAND_1028[5:0];
  _RAND_1029 = {1{`RANDOM}};
  two_complement_buffer_2_61 = _RAND_1029[5:0];
  _RAND_1030 = {1{`RANDOM}};
  two_complement_buffer_2_62 = _RAND_1030[5:0];
  _RAND_1031 = {1{`RANDOM}};
  two_complement_buffer_2_63 = _RAND_1031[5:0];
  _RAND_1032 = {1{`RANDOM}};
  multiplierReg_128 = _RAND_1032[4:0];
  _RAND_1033 = {1{`RANDOM}};
  signReg_128 = _RAND_1033[0:0];
  _RAND_1034 = {1{`RANDOM}};
  multiplierReg_129 = _RAND_1034[4:0];
  _RAND_1035 = {1{`RANDOM}};
  signReg_129 = _RAND_1035[0:0];
  _RAND_1036 = {1{`RANDOM}};
  multiplierReg_130 = _RAND_1036[4:0];
  _RAND_1037 = {1{`RANDOM}};
  signReg_130 = _RAND_1037[0:0];
  _RAND_1038 = {1{`RANDOM}};
  multiplierReg_131 = _RAND_1038[4:0];
  _RAND_1039 = {1{`RANDOM}};
  signReg_131 = _RAND_1039[0:0];
  _RAND_1040 = {1{`RANDOM}};
  multiplierReg_132 = _RAND_1040[4:0];
  _RAND_1041 = {1{`RANDOM}};
  signReg_132 = _RAND_1041[0:0];
  _RAND_1042 = {1{`RANDOM}};
  multiplierReg_133 = _RAND_1042[4:0];
  _RAND_1043 = {1{`RANDOM}};
  signReg_133 = _RAND_1043[0:0];
  _RAND_1044 = {1{`RANDOM}};
  multiplierReg_134 = _RAND_1044[4:0];
  _RAND_1045 = {1{`RANDOM}};
  signReg_134 = _RAND_1045[0:0];
  _RAND_1046 = {1{`RANDOM}};
  multiplierReg_135 = _RAND_1046[4:0];
  _RAND_1047 = {1{`RANDOM}};
  signReg_135 = _RAND_1047[0:0];
  _RAND_1048 = {1{`RANDOM}};
  multiplierReg_136 = _RAND_1048[4:0];
  _RAND_1049 = {1{`RANDOM}};
  signReg_136 = _RAND_1049[0:0];
  _RAND_1050 = {1{`RANDOM}};
  multiplierReg_137 = _RAND_1050[4:0];
  _RAND_1051 = {1{`RANDOM}};
  signReg_137 = _RAND_1051[0:0];
  _RAND_1052 = {1{`RANDOM}};
  multiplierReg_138 = _RAND_1052[4:0];
  _RAND_1053 = {1{`RANDOM}};
  signReg_138 = _RAND_1053[0:0];
  _RAND_1054 = {1{`RANDOM}};
  multiplierReg_139 = _RAND_1054[4:0];
  _RAND_1055 = {1{`RANDOM}};
  signReg_139 = _RAND_1055[0:0];
  _RAND_1056 = {1{`RANDOM}};
  multiplierReg_140 = _RAND_1056[4:0];
  _RAND_1057 = {1{`RANDOM}};
  signReg_140 = _RAND_1057[0:0];
  _RAND_1058 = {1{`RANDOM}};
  multiplierReg_141 = _RAND_1058[4:0];
  _RAND_1059 = {1{`RANDOM}};
  signReg_141 = _RAND_1059[0:0];
  _RAND_1060 = {1{`RANDOM}};
  multiplierReg_142 = _RAND_1060[4:0];
  _RAND_1061 = {1{`RANDOM}};
  signReg_142 = _RAND_1061[0:0];
  _RAND_1062 = {1{`RANDOM}};
  multiplierReg_143 = _RAND_1062[4:0];
  _RAND_1063 = {1{`RANDOM}};
  signReg_143 = _RAND_1063[0:0];
  _RAND_1064 = {1{`RANDOM}};
  multiplierReg_144 = _RAND_1064[4:0];
  _RAND_1065 = {1{`RANDOM}};
  signReg_144 = _RAND_1065[0:0];
  _RAND_1066 = {1{`RANDOM}};
  multiplierReg_145 = _RAND_1066[4:0];
  _RAND_1067 = {1{`RANDOM}};
  signReg_145 = _RAND_1067[0:0];
  _RAND_1068 = {1{`RANDOM}};
  multiplierReg_146 = _RAND_1068[4:0];
  _RAND_1069 = {1{`RANDOM}};
  signReg_146 = _RAND_1069[0:0];
  _RAND_1070 = {1{`RANDOM}};
  multiplierReg_147 = _RAND_1070[4:0];
  _RAND_1071 = {1{`RANDOM}};
  signReg_147 = _RAND_1071[0:0];
  _RAND_1072 = {1{`RANDOM}};
  multiplierReg_148 = _RAND_1072[4:0];
  _RAND_1073 = {1{`RANDOM}};
  signReg_148 = _RAND_1073[0:0];
  _RAND_1074 = {1{`RANDOM}};
  multiplierReg_149 = _RAND_1074[4:0];
  _RAND_1075 = {1{`RANDOM}};
  signReg_149 = _RAND_1075[0:0];
  _RAND_1076 = {1{`RANDOM}};
  multiplierReg_150 = _RAND_1076[4:0];
  _RAND_1077 = {1{`RANDOM}};
  signReg_150 = _RAND_1077[0:0];
  _RAND_1078 = {1{`RANDOM}};
  multiplierReg_151 = _RAND_1078[4:0];
  _RAND_1079 = {1{`RANDOM}};
  signReg_151 = _RAND_1079[0:0];
  _RAND_1080 = {1{`RANDOM}};
  multiplierReg_152 = _RAND_1080[4:0];
  _RAND_1081 = {1{`RANDOM}};
  signReg_152 = _RAND_1081[0:0];
  _RAND_1082 = {1{`RANDOM}};
  multiplierReg_153 = _RAND_1082[4:0];
  _RAND_1083 = {1{`RANDOM}};
  signReg_153 = _RAND_1083[0:0];
  _RAND_1084 = {1{`RANDOM}};
  multiplierReg_154 = _RAND_1084[4:0];
  _RAND_1085 = {1{`RANDOM}};
  signReg_154 = _RAND_1085[0:0];
  _RAND_1086 = {1{`RANDOM}};
  multiplierReg_155 = _RAND_1086[4:0];
  _RAND_1087 = {1{`RANDOM}};
  signReg_155 = _RAND_1087[0:0];
  _RAND_1088 = {1{`RANDOM}};
  multiplierReg_156 = _RAND_1088[4:0];
  _RAND_1089 = {1{`RANDOM}};
  signReg_156 = _RAND_1089[0:0];
  _RAND_1090 = {1{`RANDOM}};
  multiplierReg_157 = _RAND_1090[4:0];
  _RAND_1091 = {1{`RANDOM}};
  signReg_157 = _RAND_1091[0:0];
  _RAND_1092 = {1{`RANDOM}};
  multiplierReg_158 = _RAND_1092[4:0];
  _RAND_1093 = {1{`RANDOM}};
  signReg_158 = _RAND_1093[0:0];
  _RAND_1094 = {1{`RANDOM}};
  multiplierReg_159 = _RAND_1094[4:0];
  _RAND_1095 = {1{`RANDOM}};
  signReg_159 = _RAND_1095[0:0];
  _RAND_1096 = {1{`RANDOM}};
  multiplierReg_160 = _RAND_1096[4:0];
  _RAND_1097 = {1{`RANDOM}};
  signReg_160 = _RAND_1097[0:0];
  _RAND_1098 = {1{`RANDOM}};
  multiplierReg_161 = _RAND_1098[4:0];
  _RAND_1099 = {1{`RANDOM}};
  signReg_161 = _RAND_1099[0:0];
  _RAND_1100 = {1{`RANDOM}};
  multiplierReg_162 = _RAND_1100[4:0];
  _RAND_1101 = {1{`RANDOM}};
  signReg_162 = _RAND_1101[0:0];
  _RAND_1102 = {1{`RANDOM}};
  multiplierReg_163 = _RAND_1102[4:0];
  _RAND_1103 = {1{`RANDOM}};
  signReg_163 = _RAND_1103[0:0];
  _RAND_1104 = {1{`RANDOM}};
  multiplierReg_164 = _RAND_1104[4:0];
  _RAND_1105 = {1{`RANDOM}};
  signReg_164 = _RAND_1105[0:0];
  _RAND_1106 = {1{`RANDOM}};
  multiplierReg_165 = _RAND_1106[4:0];
  _RAND_1107 = {1{`RANDOM}};
  signReg_165 = _RAND_1107[0:0];
  _RAND_1108 = {1{`RANDOM}};
  multiplierReg_166 = _RAND_1108[4:0];
  _RAND_1109 = {1{`RANDOM}};
  signReg_166 = _RAND_1109[0:0];
  _RAND_1110 = {1{`RANDOM}};
  multiplierReg_167 = _RAND_1110[4:0];
  _RAND_1111 = {1{`RANDOM}};
  signReg_167 = _RAND_1111[0:0];
  _RAND_1112 = {1{`RANDOM}};
  multiplierReg_168 = _RAND_1112[4:0];
  _RAND_1113 = {1{`RANDOM}};
  signReg_168 = _RAND_1113[0:0];
  _RAND_1114 = {1{`RANDOM}};
  multiplierReg_169 = _RAND_1114[4:0];
  _RAND_1115 = {1{`RANDOM}};
  signReg_169 = _RAND_1115[0:0];
  _RAND_1116 = {1{`RANDOM}};
  multiplierReg_170 = _RAND_1116[4:0];
  _RAND_1117 = {1{`RANDOM}};
  signReg_170 = _RAND_1117[0:0];
  _RAND_1118 = {1{`RANDOM}};
  multiplierReg_171 = _RAND_1118[4:0];
  _RAND_1119 = {1{`RANDOM}};
  signReg_171 = _RAND_1119[0:0];
  _RAND_1120 = {1{`RANDOM}};
  multiplierReg_172 = _RAND_1120[4:0];
  _RAND_1121 = {1{`RANDOM}};
  signReg_172 = _RAND_1121[0:0];
  _RAND_1122 = {1{`RANDOM}};
  multiplierReg_173 = _RAND_1122[4:0];
  _RAND_1123 = {1{`RANDOM}};
  signReg_173 = _RAND_1123[0:0];
  _RAND_1124 = {1{`RANDOM}};
  multiplierReg_174 = _RAND_1124[4:0];
  _RAND_1125 = {1{`RANDOM}};
  signReg_174 = _RAND_1125[0:0];
  _RAND_1126 = {1{`RANDOM}};
  multiplierReg_175 = _RAND_1126[4:0];
  _RAND_1127 = {1{`RANDOM}};
  signReg_175 = _RAND_1127[0:0];
  _RAND_1128 = {1{`RANDOM}};
  multiplierReg_176 = _RAND_1128[4:0];
  _RAND_1129 = {1{`RANDOM}};
  signReg_176 = _RAND_1129[0:0];
  _RAND_1130 = {1{`RANDOM}};
  multiplierReg_177 = _RAND_1130[4:0];
  _RAND_1131 = {1{`RANDOM}};
  signReg_177 = _RAND_1131[0:0];
  _RAND_1132 = {1{`RANDOM}};
  multiplierReg_178 = _RAND_1132[4:0];
  _RAND_1133 = {1{`RANDOM}};
  signReg_178 = _RAND_1133[0:0];
  _RAND_1134 = {1{`RANDOM}};
  multiplierReg_179 = _RAND_1134[4:0];
  _RAND_1135 = {1{`RANDOM}};
  signReg_179 = _RAND_1135[0:0];
  _RAND_1136 = {1{`RANDOM}};
  multiplierReg_180 = _RAND_1136[4:0];
  _RAND_1137 = {1{`RANDOM}};
  signReg_180 = _RAND_1137[0:0];
  _RAND_1138 = {1{`RANDOM}};
  multiplierReg_181 = _RAND_1138[4:0];
  _RAND_1139 = {1{`RANDOM}};
  signReg_181 = _RAND_1139[0:0];
  _RAND_1140 = {1{`RANDOM}};
  multiplierReg_182 = _RAND_1140[4:0];
  _RAND_1141 = {1{`RANDOM}};
  signReg_182 = _RAND_1141[0:0];
  _RAND_1142 = {1{`RANDOM}};
  multiplierReg_183 = _RAND_1142[4:0];
  _RAND_1143 = {1{`RANDOM}};
  signReg_183 = _RAND_1143[0:0];
  _RAND_1144 = {1{`RANDOM}};
  multiplierReg_184 = _RAND_1144[4:0];
  _RAND_1145 = {1{`RANDOM}};
  signReg_184 = _RAND_1145[0:0];
  _RAND_1146 = {1{`RANDOM}};
  multiplierReg_185 = _RAND_1146[4:0];
  _RAND_1147 = {1{`RANDOM}};
  signReg_185 = _RAND_1147[0:0];
  _RAND_1148 = {1{`RANDOM}};
  multiplierReg_186 = _RAND_1148[4:0];
  _RAND_1149 = {1{`RANDOM}};
  signReg_186 = _RAND_1149[0:0];
  _RAND_1150 = {1{`RANDOM}};
  multiplierReg_187 = _RAND_1150[4:0];
  _RAND_1151 = {1{`RANDOM}};
  signReg_187 = _RAND_1151[0:0];
  _RAND_1152 = {1{`RANDOM}};
  multiplierReg_188 = _RAND_1152[4:0];
  _RAND_1153 = {1{`RANDOM}};
  signReg_188 = _RAND_1153[0:0];
  _RAND_1154 = {1{`RANDOM}};
  multiplierReg_189 = _RAND_1154[4:0];
  _RAND_1155 = {1{`RANDOM}};
  signReg_189 = _RAND_1155[0:0];
  _RAND_1156 = {1{`RANDOM}};
  multiplierReg_190 = _RAND_1156[4:0];
  _RAND_1157 = {1{`RANDOM}};
  signReg_190 = _RAND_1157[0:0];
  _RAND_1158 = {1{`RANDOM}};
  multiplierReg_191 = _RAND_1158[4:0];
  _RAND_1159 = {1{`RANDOM}};
  signReg_191 = _RAND_1159[0:0];
  _RAND_1160 = {1{`RANDOM}};
  dotProductRegs_3_0 = _RAND_1160[4:0];
  _RAND_1161 = {1{`RANDOM}};
  dotProductRegs_3_1 = _RAND_1161[4:0];
  _RAND_1162 = {1{`RANDOM}};
  dotProductRegs_3_2 = _RAND_1162[4:0];
  _RAND_1163 = {1{`RANDOM}};
  dotProductRegs_3_3 = _RAND_1163[4:0];
  _RAND_1164 = {1{`RANDOM}};
  dotProductRegs_3_4 = _RAND_1164[4:0];
  _RAND_1165 = {1{`RANDOM}};
  dotProductRegs_3_5 = _RAND_1165[4:0];
  _RAND_1166 = {1{`RANDOM}};
  dotProductRegs_3_6 = _RAND_1166[4:0];
  _RAND_1167 = {1{`RANDOM}};
  dotProductRegs_3_7 = _RAND_1167[4:0];
  _RAND_1168 = {1{`RANDOM}};
  dotProductRegs_3_8 = _RAND_1168[4:0];
  _RAND_1169 = {1{`RANDOM}};
  dotProductRegs_3_9 = _RAND_1169[4:0];
  _RAND_1170 = {1{`RANDOM}};
  dotProductRegs_3_10 = _RAND_1170[4:0];
  _RAND_1171 = {1{`RANDOM}};
  dotProductRegs_3_11 = _RAND_1171[4:0];
  _RAND_1172 = {1{`RANDOM}};
  dotProductRegs_3_12 = _RAND_1172[4:0];
  _RAND_1173 = {1{`RANDOM}};
  dotProductRegs_3_13 = _RAND_1173[4:0];
  _RAND_1174 = {1{`RANDOM}};
  dotProductRegs_3_14 = _RAND_1174[4:0];
  _RAND_1175 = {1{`RANDOM}};
  dotProductRegs_3_15 = _RAND_1175[4:0];
  _RAND_1176 = {1{`RANDOM}};
  dotProductRegs_3_16 = _RAND_1176[4:0];
  _RAND_1177 = {1{`RANDOM}};
  dotProductRegs_3_17 = _RAND_1177[4:0];
  _RAND_1178 = {1{`RANDOM}};
  dotProductRegs_3_18 = _RAND_1178[4:0];
  _RAND_1179 = {1{`RANDOM}};
  dotProductRegs_3_19 = _RAND_1179[4:0];
  _RAND_1180 = {1{`RANDOM}};
  dotProductRegs_3_20 = _RAND_1180[4:0];
  _RAND_1181 = {1{`RANDOM}};
  dotProductRegs_3_21 = _RAND_1181[4:0];
  _RAND_1182 = {1{`RANDOM}};
  dotProductRegs_3_22 = _RAND_1182[4:0];
  _RAND_1183 = {1{`RANDOM}};
  dotProductRegs_3_23 = _RAND_1183[4:0];
  _RAND_1184 = {1{`RANDOM}};
  dotProductRegs_3_24 = _RAND_1184[4:0];
  _RAND_1185 = {1{`RANDOM}};
  dotProductRegs_3_25 = _RAND_1185[4:0];
  _RAND_1186 = {1{`RANDOM}};
  dotProductRegs_3_26 = _RAND_1186[4:0];
  _RAND_1187 = {1{`RANDOM}};
  dotProductRegs_3_27 = _RAND_1187[4:0];
  _RAND_1188 = {1{`RANDOM}};
  dotProductRegs_3_28 = _RAND_1188[4:0];
  _RAND_1189 = {1{`RANDOM}};
  dotProductRegs_3_29 = _RAND_1189[4:0];
  _RAND_1190 = {1{`RANDOM}};
  dotProductRegs_3_30 = _RAND_1190[4:0];
  _RAND_1191 = {1{`RANDOM}};
  dotProductRegs_3_31 = _RAND_1191[4:0];
  _RAND_1192 = {1{`RANDOM}};
  dotProductRegs_3_32 = _RAND_1192[4:0];
  _RAND_1193 = {1{`RANDOM}};
  dotProductRegs_3_33 = _RAND_1193[4:0];
  _RAND_1194 = {1{`RANDOM}};
  dotProductRegs_3_34 = _RAND_1194[4:0];
  _RAND_1195 = {1{`RANDOM}};
  dotProductRegs_3_35 = _RAND_1195[4:0];
  _RAND_1196 = {1{`RANDOM}};
  dotProductRegs_3_36 = _RAND_1196[4:0];
  _RAND_1197 = {1{`RANDOM}};
  dotProductRegs_3_37 = _RAND_1197[4:0];
  _RAND_1198 = {1{`RANDOM}};
  dotProductRegs_3_38 = _RAND_1198[4:0];
  _RAND_1199 = {1{`RANDOM}};
  dotProductRegs_3_39 = _RAND_1199[4:0];
  _RAND_1200 = {1{`RANDOM}};
  dotProductRegs_3_40 = _RAND_1200[4:0];
  _RAND_1201 = {1{`RANDOM}};
  dotProductRegs_3_41 = _RAND_1201[4:0];
  _RAND_1202 = {1{`RANDOM}};
  dotProductRegs_3_42 = _RAND_1202[4:0];
  _RAND_1203 = {1{`RANDOM}};
  dotProductRegs_3_43 = _RAND_1203[4:0];
  _RAND_1204 = {1{`RANDOM}};
  dotProductRegs_3_44 = _RAND_1204[4:0];
  _RAND_1205 = {1{`RANDOM}};
  dotProductRegs_3_45 = _RAND_1205[4:0];
  _RAND_1206 = {1{`RANDOM}};
  dotProductRegs_3_46 = _RAND_1206[4:0];
  _RAND_1207 = {1{`RANDOM}};
  dotProductRegs_3_47 = _RAND_1207[4:0];
  _RAND_1208 = {1{`RANDOM}};
  dotProductRegs_3_48 = _RAND_1208[4:0];
  _RAND_1209 = {1{`RANDOM}};
  dotProductRegs_3_49 = _RAND_1209[4:0];
  _RAND_1210 = {1{`RANDOM}};
  dotProductRegs_3_50 = _RAND_1210[4:0];
  _RAND_1211 = {1{`RANDOM}};
  dotProductRegs_3_51 = _RAND_1211[4:0];
  _RAND_1212 = {1{`RANDOM}};
  dotProductRegs_3_52 = _RAND_1212[4:0];
  _RAND_1213 = {1{`RANDOM}};
  dotProductRegs_3_53 = _RAND_1213[4:0];
  _RAND_1214 = {1{`RANDOM}};
  dotProductRegs_3_54 = _RAND_1214[4:0];
  _RAND_1215 = {1{`RANDOM}};
  dotProductRegs_3_55 = _RAND_1215[4:0];
  _RAND_1216 = {1{`RANDOM}};
  dotProductRegs_3_56 = _RAND_1216[4:0];
  _RAND_1217 = {1{`RANDOM}};
  dotProductRegs_3_57 = _RAND_1217[4:0];
  _RAND_1218 = {1{`RANDOM}};
  dotProductRegs_3_58 = _RAND_1218[4:0];
  _RAND_1219 = {1{`RANDOM}};
  dotProductRegs_3_59 = _RAND_1219[4:0];
  _RAND_1220 = {1{`RANDOM}};
  dotProductRegs_3_60 = _RAND_1220[4:0];
  _RAND_1221 = {1{`RANDOM}};
  dotProductRegs_3_61 = _RAND_1221[4:0];
  _RAND_1222 = {1{`RANDOM}};
  dotProductRegs_3_62 = _RAND_1222[4:0];
  _RAND_1223 = {1{`RANDOM}};
  dotProductRegs_3_63 = _RAND_1223[4:0];
  _RAND_1224 = {1{`RANDOM}};
  signs_3_0 = _RAND_1224[0:0];
  _RAND_1225 = {1{`RANDOM}};
  signs_3_1 = _RAND_1225[0:0];
  _RAND_1226 = {1{`RANDOM}};
  signs_3_2 = _RAND_1226[0:0];
  _RAND_1227 = {1{`RANDOM}};
  signs_3_3 = _RAND_1227[0:0];
  _RAND_1228 = {1{`RANDOM}};
  signs_3_4 = _RAND_1228[0:0];
  _RAND_1229 = {1{`RANDOM}};
  signs_3_5 = _RAND_1229[0:0];
  _RAND_1230 = {1{`RANDOM}};
  signs_3_6 = _RAND_1230[0:0];
  _RAND_1231 = {1{`RANDOM}};
  signs_3_7 = _RAND_1231[0:0];
  _RAND_1232 = {1{`RANDOM}};
  signs_3_8 = _RAND_1232[0:0];
  _RAND_1233 = {1{`RANDOM}};
  signs_3_9 = _RAND_1233[0:0];
  _RAND_1234 = {1{`RANDOM}};
  signs_3_10 = _RAND_1234[0:0];
  _RAND_1235 = {1{`RANDOM}};
  signs_3_11 = _RAND_1235[0:0];
  _RAND_1236 = {1{`RANDOM}};
  signs_3_12 = _RAND_1236[0:0];
  _RAND_1237 = {1{`RANDOM}};
  signs_3_13 = _RAND_1237[0:0];
  _RAND_1238 = {1{`RANDOM}};
  signs_3_14 = _RAND_1238[0:0];
  _RAND_1239 = {1{`RANDOM}};
  signs_3_15 = _RAND_1239[0:0];
  _RAND_1240 = {1{`RANDOM}};
  signs_3_16 = _RAND_1240[0:0];
  _RAND_1241 = {1{`RANDOM}};
  signs_3_17 = _RAND_1241[0:0];
  _RAND_1242 = {1{`RANDOM}};
  signs_3_18 = _RAND_1242[0:0];
  _RAND_1243 = {1{`RANDOM}};
  signs_3_19 = _RAND_1243[0:0];
  _RAND_1244 = {1{`RANDOM}};
  signs_3_20 = _RAND_1244[0:0];
  _RAND_1245 = {1{`RANDOM}};
  signs_3_21 = _RAND_1245[0:0];
  _RAND_1246 = {1{`RANDOM}};
  signs_3_22 = _RAND_1246[0:0];
  _RAND_1247 = {1{`RANDOM}};
  signs_3_23 = _RAND_1247[0:0];
  _RAND_1248 = {1{`RANDOM}};
  signs_3_24 = _RAND_1248[0:0];
  _RAND_1249 = {1{`RANDOM}};
  signs_3_25 = _RAND_1249[0:0];
  _RAND_1250 = {1{`RANDOM}};
  signs_3_26 = _RAND_1250[0:0];
  _RAND_1251 = {1{`RANDOM}};
  signs_3_27 = _RAND_1251[0:0];
  _RAND_1252 = {1{`RANDOM}};
  signs_3_28 = _RAND_1252[0:0];
  _RAND_1253 = {1{`RANDOM}};
  signs_3_29 = _RAND_1253[0:0];
  _RAND_1254 = {1{`RANDOM}};
  signs_3_30 = _RAND_1254[0:0];
  _RAND_1255 = {1{`RANDOM}};
  signs_3_31 = _RAND_1255[0:0];
  _RAND_1256 = {1{`RANDOM}};
  signs_3_32 = _RAND_1256[0:0];
  _RAND_1257 = {1{`RANDOM}};
  signs_3_33 = _RAND_1257[0:0];
  _RAND_1258 = {1{`RANDOM}};
  signs_3_34 = _RAND_1258[0:0];
  _RAND_1259 = {1{`RANDOM}};
  signs_3_35 = _RAND_1259[0:0];
  _RAND_1260 = {1{`RANDOM}};
  signs_3_36 = _RAND_1260[0:0];
  _RAND_1261 = {1{`RANDOM}};
  signs_3_37 = _RAND_1261[0:0];
  _RAND_1262 = {1{`RANDOM}};
  signs_3_38 = _RAND_1262[0:0];
  _RAND_1263 = {1{`RANDOM}};
  signs_3_39 = _RAND_1263[0:0];
  _RAND_1264 = {1{`RANDOM}};
  signs_3_40 = _RAND_1264[0:0];
  _RAND_1265 = {1{`RANDOM}};
  signs_3_41 = _RAND_1265[0:0];
  _RAND_1266 = {1{`RANDOM}};
  signs_3_42 = _RAND_1266[0:0];
  _RAND_1267 = {1{`RANDOM}};
  signs_3_43 = _RAND_1267[0:0];
  _RAND_1268 = {1{`RANDOM}};
  signs_3_44 = _RAND_1268[0:0];
  _RAND_1269 = {1{`RANDOM}};
  signs_3_45 = _RAND_1269[0:0];
  _RAND_1270 = {1{`RANDOM}};
  signs_3_46 = _RAND_1270[0:0];
  _RAND_1271 = {1{`RANDOM}};
  signs_3_47 = _RAND_1271[0:0];
  _RAND_1272 = {1{`RANDOM}};
  signs_3_48 = _RAND_1272[0:0];
  _RAND_1273 = {1{`RANDOM}};
  signs_3_49 = _RAND_1273[0:0];
  _RAND_1274 = {1{`RANDOM}};
  signs_3_50 = _RAND_1274[0:0];
  _RAND_1275 = {1{`RANDOM}};
  signs_3_51 = _RAND_1275[0:0];
  _RAND_1276 = {1{`RANDOM}};
  signs_3_52 = _RAND_1276[0:0];
  _RAND_1277 = {1{`RANDOM}};
  signs_3_53 = _RAND_1277[0:0];
  _RAND_1278 = {1{`RANDOM}};
  signs_3_54 = _RAND_1278[0:0];
  _RAND_1279 = {1{`RANDOM}};
  signs_3_55 = _RAND_1279[0:0];
  _RAND_1280 = {1{`RANDOM}};
  signs_3_56 = _RAND_1280[0:0];
  _RAND_1281 = {1{`RANDOM}};
  signs_3_57 = _RAND_1281[0:0];
  _RAND_1282 = {1{`RANDOM}};
  signs_3_58 = _RAND_1282[0:0];
  _RAND_1283 = {1{`RANDOM}};
  signs_3_59 = _RAND_1283[0:0];
  _RAND_1284 = {1{`RANDOM}};
  signs_3_60 = _RAND_1284[0:0];
  _RAND_1285 = {1{`RANDOM}};
  signs_3_61 = _RAND_1285[0:0];
  _RAND_1286 = {1{`RANDOM}};
  signs_3_62 = _RAND_1286[0:0];
  _RAND_1287 = {1{`RANDOM}};
  signs_3_63 = _RAND_1287[0:0];
  _RAND_1288 = {1{`RANDOM}};
  two_complement_3_0 = _RAND_1288[5:0];
  _RAND_1289 = {1{`RANDOM}};
  two_complement_3_1 = _RAND_1289[5:0];
  _RAND_1290 = {1{`RANDOM}};
  two_complement_3_2 = _RAND_1290[5:0];
  _RAND_1291 = {1{`RANDOM}};
  two_complement_3_3 = _RAND_1291[5:0];
  _RAND_1292 = {1{`RANDOM}};
  two_complement_3_4 = _RAND_1292[5:0];
  _RAND_1293 = {1{`RANDOM}};
  two_complement_3_5 = _RAND_1293[5:0];
  _RAND_1294 = {1{`RANDOM}};
  two_complement_3_6 = _RAND_1294[5:0];
  _RAND_1295 = {1{`RANDOM}};
  two_complement_3_7 = _RAND_1295[5:0];
  _RAND_1296 = {1{`RANDOM}};
  two_complement_3_8 = _RAND_1296[5:0];
  _RAND_1297 = {1{`RANDOM}};
  two_complement_3_9 = _RAND_1297[5:0];
  _RAND_1298 = {1{`RANDOM}};
  two_complement_3_10 = _RAND_1298[5:0];
  _RAND_1299 = {1{`RANDOM}};
  two_complement_3_11 = _RAND_1299[5:0];
  _RAND_1300 = {1{`RANDOM}};
  two_complement_3_12 = _RAND_1300[5:0];
  _RAND_1301 = {1{`RANDOM}};
  two_complement_3_13 = _RAND_1301[5:0];
  _RAND_1302 = {1{`RANDOM}};
  two_complement_3_14 = _RAND_1302[5:0];
  _RAND_1303 = {1{`RANDOM}};
  two_complement_3_15 = _RAND_1303[5:0];
  _RAND_1304 = {1{`RANDOM}};
  two_complement_3_16 = _RAND_1304[5:0];
  _RAND_1305 = {1{`RANDOM}};
  two_complement_3_17 = _RAND_1305[5:0];
  _RAND_1306 = {1{`RANDOM}};
  two_complement_3_18 = _RAND_1306[5:0];
  _RAND_1307 = {1{`RANDOM}};
  two_complement_3_19 = _RAND_1307[5:0];
  _RAND_1308 = {1{`RANDOM}};
  two_complement_3_20 = _RAND_1308[5:0];
  _RAND_1309 = {1{`RANDOM}};
  two_complement_3_21 = _RAND_1309[5:0];
  _RAND_1310 = {1{`RANDOM}};
  two_complement_3_22 = _RAND_1310[5:0];
  _RAND_1311 = {1{`RANDOM}};
  two_complement_3_23 = _RAND_1311[5:0];
  _RAND_1312 = {1{`RANDOM}};
  two_complement_3_24 = _RAND_1312[5:0];
  _RAND_1313 = {1{`RANDOM}};
  two_complement_3_25 = _RAND_1313[5:0];
  _RAND_1314 = {1{`RANDOM}};
  two_complement_3_26 = _RAND_1314[5:0];
  _RAND_1315 = {1{`RANDOM}};
  two_complement_3_27 = _RAND_1315[5:0];
  _RAND_1316 = {1{`RANDOM}};
  two_complement_3_28 = _RAND_1316[5:0];
  _RAND_1317 = {1{`RANDOM}};
  two_complement_3_29 = _RAND_1317[5:0];
  _RAND_1318 = {1{`RANDOM}};
  two_complement_3_30 = _RAND_1318[5:0];
  _RAND_1319 = {1{`RANDOM}};
  two_complement_3_31 = _RAND_1319[5:0];
  _RAND_1320 = {1{`RANDOM}};
  two_complement_3_32 = _RAND_1320[5:0];
  _RAND_1321 = {1{`RANDOM}};
  two_complement_3_33 = _RAND_1321[5:0];
  _RAND_1322 = {1{`RANDOM}};
  two_complement_3_34 = _RAND_1322[5:0];
  _RAND_1323 = {1{`RANDOM}};
  two_complement_3_35 = _RAND_1323[5:0];
  _RAND_1324 = {1{`RANDOM}};
  two_complement_3_36 = _RAND_1324[5:0];
  _RAND_1325 = {1{`RANDOM}};
  two_complement_3_37 = _RAND_1325[5:0];
  _RAND_1326 = {1{`RANDOM}};
  two_complement_3_38 = _RAND_1326[5:0];
  _RAND_1327 = {1{`RANDOM}};
  two_complement_3_39 = _RAND_1327[5:0];
  _RAND_1328 = {1{`RANDOM}};
  two_complement_3_40 = _RAND_1328[5:0];
  _RAND_1329 = {1{`RANDOM}};
  two_complement_3_41 = _RAND_1329[5:0];
  _RAND_1330 = {1{`RANDOM}};
  two_complement_3_42 = _RAND_1330[5:0];
  _RAND_1331 = {1{`RANDOM}};
  two_complement_3_43 = _RAND_1331[5:0];
  _RAND_1332 = {1{`RANDOM}};
  two_complement_3_44 = _RAND_1332[5:0];
  _RAND_1333 = {1{`RANDOM}};
  two_complement_3_45 = _RAND_1333[5:0];
  _RAND_1334 = {1{`RANDOM}};
  two_complement_3_46 = _RAND_1334[5:0];
  _RAND_1335 = {1{`RANDOM}};
  two_complement_3_47 = _RAND_1335[5:0];
  _RAND_1336 = {1{`RANDOM}};
  two_complement_3_48 = _RAND_1336[5:0];
  _RAND_1337 = {1{`RANDOM}};
  two_complement_3_49 = _RAND_1337[5:0];
  _RAND_1338 = {1{`RANDOM}};
  two_complement_3_50 = _RAND_1338[5:0];
  _RAND_1339 = {1{`RANDOM}};
  two_complement_3_51 = _RAND_1339[5:0];
  _RAND_1340 = {1{`RANDOM}};
  two_complement_3_52 = _RAND_1340[5:0];
  _RAND_1341 = {1{`RANDOM}};
  two_complement_3_53 = _RAND_1341[5:0];
  _RAND_1342 = {1{`RANDOM}};
  two_complement_3_54 = _RAND_1342[5:0];
  _RAND_1343 = {1{`RANDOM}};
  two_complement_3_55 = _RAND_1343[5:0];
  _RAND_1344 = {1{`RANDOM}};
  two_complement_3_56 = _RAND_1344[5:0];
  _RAND_1345 = {1{`RANDOM}};
  two_complement_3_57 = _RAND_1345[5:0];
  _RAND_1346 = {1{`RANDOM}};
  two_complement_3_58 = _RAND_1346[5:0];
  _RAND_1347 = {1{`RANDOM}};
  two_complement_3_59 = _RAND_1347[5:0];
  _RAND_1348 = {1{`RANDOM}};
  two_complement_3_60 = _RAND_1348[5:0];
  _RAND_1349 = {1{`RANDOM}};
  two_complement_3_61 = _RAND_1349[5:0];
  _RAND_1350 = {1{`RANDOM}};
  two_complement_3_62 = _RAND_1350[5:0];
  _RAND_1351 = {1{`RANDOM}};
  two_complement_3_63 = _RAND_1351[5:0];
  _RAND_1352 = {1{`RANDOM}};
  two_complement_buffer_3_0 = _RAND_1352[5:0];
  _RAND_1353 = {1{`RANDOM}};
  two_complement_buffer_3_1 = _RAND_1353[5:0];
  _RAND_1354 = {1{`RANDOM}};
  two_complement_buffer_3_2 = _RAND_1354[5:0];
  _RAND_1355 = {1{`RANDOM}};
  two_complement_buffer_3_3 = _RAND_1355[5:0];
  _RAND_1356 = {1{`RANDOM}};
  two_complement_buffer_3_4 = _RAND_1356[5:0];
  _RAND_1357 = {1{`RANDOM}};
  two_complement_buffer_3_5 = _RAND_1357[5:0];
  _RAND_1358 = {1{`RANDOM}};
  two_complement_buffer_3_6 = _RAND_1358[5:0];
  _RAND_1359 = {1{`RANDOM}};
  two_complement_buffer_3_7 = _RAND_1359[5:0];
  _RAND_1360 = {1{`RANDOM}};
  two_complement_buffer_3_8 = _RAND_1360[5:0];
  _RAND_1361 = {1{`RANDOM}};
  two_complement_buffer_3_9 = _RAND_1361[5:0];
  _RAND_1362 = {1{`RANDOM}};
  two_complement_buffer_3_10 = _RAND_1362[5:0];
  _RAND_1363 = {1{`RANDOM}};
  two_complement_buffer_3_11 = _RAND_1363[5:0];
  _RAND_1364 = {1{`RANDOM}};
  two_complement_buffer_3_12 = _RAND_1364[5:0];
  _RAND_1365 = {1{`RANDOM}};
  two_complement_buffer_3_13 = _RAND_1365[5:0];
  _RAND_1366 = {1{`RANDOM}};
  two_complement_buffer_3_14 = _RAND_1366[5:0];
  _RAND_1367 = {1{`RANDOM}};
  two_complement_buffer_3_15 = _RAND_1367[5:0];
  _RAND_1368 = {1{`RANDOM}};
  two_complement_buffer_3_16 = _RAND_1368[5:0];
  _RAND_1369 = {1{`RANDOM}};
  two_complement_buffer_3_17 = _RAND_1369[5:0];
  _RAND_1370 = {1{`RANDOM}};
  two_complement_buffer_3_18 = _RAND_1370[5:0];
  _RAND_1371 = {1{`RANDOM}};
  two_complement_buffer_3_19 = _RAND_1371[5:0];
  _RAND_1372 = {1{`RANDOM}};
  two_complement_buffer_3_20 = _RAND_1372[5:0];
  _RAND_1373 = {1{`RANDOM}};
  two_complement_buffer_3_21 = _RAND_1373[5:0];
  _RAND_1374 = {1{`RANDOM}};
  two_complement_buffer_3_22 = _RAND_1374[5:0];
  _RAND_1375 = {1{`RANDOM}};
  two_complement_buffer_3_23 = _RAND_1375[5:0];
  _RAND_1376 = {1{`RANDOM}};
  two_complement_buffer_3_24 = _RAND_1376[5:0];
  _RAND_1377 = {1{`RANDOM}};
  two_complement_buffer_3_25 = _RAND_1377[5:0];
  _RAND_1378 = {1{`RANDOM}};
  two_complement_buffer_3_26 = _RAND_1378[5:0];
  _RAND_1379 = {1{`RANDOM}};
  two_complement_buffer_3_27 = _RAND_1379[5:0];
  _RAND_1380 = {1{`RANDOM}};
  two_complement_buffer_3_28 = _RAND_1380[5:0];
  _RAND_1381 = {1{`RANDOM}};
  two_complement_buffer_3_29 = _RAND_1381[5:0];
  _RAND_1382 = {1{`RANDOM}};
  two_complement_buffer_3_30 = _RAND_1382[5:0];
  _RAND_1383 = {1{`RANDOM}};
  two_complement_buffer_3_31 = _RAND_1383[5:0];
  _RAND_1384 = {1{`RANDOM}};
  two_complement_buffer_3_32 = _RAND_1384[5:0];
  _RAND_1385 = {1{`RANDOM}};
  two_complement_buffer_3_33 = _RAND_1385[5:0];
  _RAND_1386 = {1{`RANDOM}};
  two_complement_buffer_3_34 = _RAND_1386[5:0];
  _RAND_1387 = {1{`RANDOM}};
  two_complement_buffer_3_35 = _RAND_1387[5:0];
  _RAND_1388 = {1{`RANDOM}};
  two_complement_buffer_3_36 = _RAND_1388[5:0];
  _RAND_1389 = {1{`RANDOM}};
  two_complement_buffer_3_37 = _RAND_1389[5:0];
  _RAND_1390 = {1{`RANDOM}};
  two_complement_buffer_3_38 = _RAND_1390[5:0];
  _RAND_1391 = {1{`RANDOM}};
  two_complement_buffer_3_39 = _RAND_1391[5:0];
  _RAND_1392 = {1{`RANDOM}};
  two_complement_buffer_3_40 = _RAND_1392[5:0];
  _RAND_1393 = {1{`RANDOM}};
  two_complement_buffer_3_41 = _RAND_1393[5:0];
  _RAND_1394 = {1{`RANDOM}};
  two_complement_buffer_3_42 = _RAND_1394[5:0];
  _RAND_1395 = {1{`RANDOM}};
  two_complement_buffer_3_43 = _RAND_1395[5:0];
  _RAND_1396 = {1{`RANDOM}};
  two_complement_buffer_3_44 = _RAND_1396[5:0];
  _RAND_1397 = {1{`RANDOM}};
  two_complement_buffer_3_45 = _RAND_1397[5:0];
  _RAND_1398 = {1{`RANDOM}};
  two_complement_buffer_3_46 = _RAND_1398[5:0];
  _RAND_1399 = {1{`RANDOM}};
  two_complement_buffer_3_47 = _RAND_1399[5:0];
  _RAND_1400 = {1{`RANDOM}};
  two_complement_buffer_3_48 = _RAND_1400[5:0];
  _RAND_1401 = {1{`RANDOM}};
  two_complement_buffer_3_49 = _RAND_1401[5:0];
  _RAND_1402 = {1{`RANDOM}};
  two_complement_buffer_3_50 = _RAND_1402[5:0];
  _RAND_1403 = {1{`RANDOM}};
  two_complement_buffer_3_51 = _RAND_1403[5:0];
  _RAND_1404 = {1{`RANDOM}};
  two_complement_buffer_3_52 = _RAND_1404[5:0];
  _RAND_1405 = {1{`RANDOM}};
  two_complement_buffer_3_53 = _RAND_1405[5:0];
  _RAND_1406 = {1{`RANDOM}};
  two_complement_buffer_3_54 = _RAND_1406[5:0];
  _RAND_1407 = {1{`RANDOM}};
  two_complement_buffer_3_55 = _RAND_1407[5:0];
  _RAND_1408 = {1{`RANDOM}};
  two_complement_buffer_3_56 = _RAND_1408[5:0];
  _RAND_1409 = {1{`RANDOM}};
  two_complement_buffer_3_57 = _RAND_1409[5:0];
  _RAND_1410 = {1{`RANDOM}};
  two_complement_buffer_3_58 = _RAND_1410[5:0];
  _RAND_1411 = {1{`RANDOM}};
  two_complement_buffer_3_59 = _RAND_1411[5:0];
  _RAND_1412 = {1{`RANDOM}};
  two_complement_buffer_3_60 = _RAND_1412[5:0];
  _RAND_1413 = {1{`RANDOM}};
  two_complement_buffer_3_61 = _RAND_1413[5:0];
  _RAND_1414 = {1{`RANDOM}};
  two_complement_buffer_3_62 = _RAND_1414[5:0];
  _RAND_1415 = {1{`RANDOM}};
  two_complement_buffer_3_63 = _RAND_1415[5:0];
  _RAND_1416 = {1{`RANDOM}};
  multiplierReg_192 = _RAND_1416[4:0];
  _RAND_1417 = {1{`RANDOM}};
  signReg_192 = _RAND_1417[0:0];
  _RAND_1418 = {1{`RANDOM}};
  multiplierReg_193 = _RAND_1418[4:0];
  _RAND_1419 = {1{`RANDOM}};
  signReg_193 = _RAND_1419[0:0];
  _RAND_1420 = {1{`RANDOM}};
  multiplierReg_194 = _RAND_1420[4:0];
  _RAND_1421 = {1{`RANDOM}};
  signReg_194 = _RAND_1421[0:0];
  _RAND_1422 = {1{`RANDOM}};
  multiplierReg_195 = _RAND_1422[4:0];
  _RAND_1423 = {1{`RANDOM}};
  signReg_195 = _RAND_1423[0:0];
  _RAND_1424 = {1{`RANDOM}};
  multiplierReg_196 = _RAND_1424[4:0];
  _RAND_1425 = {1{`RANDOM}};
  signReg_196 = _RAND_1425[0:0];
  _RAND_1426 = {1{`RANDOM}};
  multiplierReg_197 = _RAND_1426[4:0];
  _RAND_1427 = {1{`RANDOM}};
  signReg_197 = _RAND_1427[0:0];
  _RAND_1428 = {1{`RANDOM}};
  multiplierReg_198 = _RAND_1428[4:0];
  _RAND_1429 = {1{`RANDOM}};
  signReg_198 = _RAND_1429[0:0];
  _RAND_1430 = {1{`RANDOM}};
  multiplierReg_199 = _RAND_1430[4:0];
  _RAND_1431 = {1{`RANDOM}};
  signReg_199 = _RAND_1431[0:0];
  _RAND_1432 = {1{`RANDOM}};
  multiplierReg_200 = _RAND_1432[4:0];
  _RAND_1433 = {1{`RANDOM}};
  signReg_200 = _RAND_1433[0:0];
  _RAND_1434 = {1{`RANDOM}};
  multiplierReg_201 = _RAND_1434[4:0];
  _RAND_1435 = {1{`RANDOM}};
  signReg_201 = _RAND_1435[0:0];
  _RAND_1436 = {1{`RANDOM}};
  multiplierReg_202 = _RAND_1436[4:0];
  _RAND_1437 = {1{`RANDOM}};
  signReg_202 = _RAND_1437[0:0];
  _RAND_1438 = {1{`RANDOM}};
  multiplierReg_203 = _RAND_1438[4:0];
  _RAND_1439 = {1{`RANDOM}};
  signReg_203 = _RAND_1439[0:0];
  _RAND_1440 = {1{`RANDOM}};
  multiplierReg_204 = _RAND_1440[4:0];
  _RAND_1441 = {1{`RANDOM}};
  signReg_204 = _RAND_1441[0:0];
  _RAND_1442 = {1{`RANDOM}};
  multiplierReg_205 = _RAND_1442[4:0];
  _RAND_1443 = {1{`RANDOM}};
  signReg_205 = _RAND_1443[0:0];
  _RAND_1444 = {1{`RANDOM}};
  multiplierReg_206 = _RAND_1444[4:0];
  _RAND_1445 = {1{`RANDOM}};
  signReg_206 = _RAND_1445[0:0];
  _RAND_1446 = {1{`RANDOM}};
  multiplierReg_207 = _RAND_1446[4:0];
  _RAND_1447 = {1{`RANDOM}};
  signReg_207 = _RAND_1447[0:0];
  _RAND_1448 = {1{`RANDOM}};
  multiplierReg_208 = _RAND_1448[4:0];
  _RAND_1449 = {1{`RANDOM}};
  signReg_208 = _RAND_1449[0:0];
  _RAND_1450 = {1{`RANDOM}};
  multiplierReg_209 = _RAND_1450[4:0];
  _RAND_1451 = {1{`RANDOM}};
  signReg_209 = _RAND_1451[0:0];
  _RAND_1452 = {1{`RANDOM}};
  multiplierReg_210 = _RAND_1452[4:0];
  _RAND_1453 = {1{`RANDOM}};
  signReg_210 = _RAND_1453[0:0];
  _RAND_1454 = {1{`RANDOM}};
  multiplierReg_211 = _RAND_1454[4:0];
  _RAND_1455 = {1{`RANDOM}};
  signReg_211 = _RAND_1455[0:0];
  _RAND_1456 = {1{`RANDOM}};
  multiplierReg_212 = _RAND_1456[4:0];
  _RAND_1457 = {1{`RANDOM}};
  signReg_212 = _RAND_1457[0:0];
  _RAND_1458 = {1{`RANDOM}};
  multiplierReg_213 = _RAND_1458[4:0];
  _RAND_1459 = {1{`RANDOM}};
  signReg_213 = _RAND_1459[0:0];
  _RAND_1460 = {1{`RANDOM}};
  multiplierReg_214 = _RAND_1460[4:0];
  _RAND_1461 = {1{`RANDOM}};
  signReg_214 = _RAND_1461[0:0];
  _RAND_1462 = {1{`RANDOM}};
  multiplierReg_215 = _RAND_1462[4:0];
  _RAND_1463 = {1{`RANDOM}};
  signReg_215 = _RAND_1463[0:0];
  _RAND_1464 = {1{`RANDOM}};
  multiplierReg_216 = _RAND_1464[4:0];
  _RAND_1465 = {1{`RANDOM}};
  signReg_216 = _RAND_1465[0:0];
  _RAND_1466 = {1{`RANDOM}};
  multiplierReg_217 = _RAND_1466[4:0];
  _RAND_1467 = {1{`RANDOM}};
  signReg_217 = _RAND_1467[0:0];
  _RAND_1468 = {1{`RANDOM}};
  multiplierReg_218 = _RAND_1468[4:0];
  _RAND_1469 = {1{`RANDOM}};
  signReg_218 = _RAND_1469[0:0];
  _RAND_1470 = {1{`RANDOM}};
  multiplierReg_219 = _RAND_1470[4:0];
  _RAND_1471 = {1{`RANDOM}};
  signReg_219 = _RAND_1471[0:0];
  _RAND_1472 = {1{`RANDOM}};
  multiplierReg_220 = _RAND_1472[4:0];
  _RAND_1473 = {1{`RANDOM}};
  signReg_220 = _RAND_1473[0:0];
  _RAND_1474 = {1{`RANDOM}};
  multiplierReg_221 = _RAND_1474[4:0];
  _RAND_1475 = {1{`RANDOM}};
  signReg_221 = _RAND_1475[0:0];
  _RAND_1476 = {1{`RANDOM}};
  multiplierReg_222 = _RAND_1476[4:0];
  _RAND_1477 = {1{`RANDOM}};
  signReg_222 = _RAND_1477[0:0];
  _RAND_1478 = {1{`RANDOM}};
  multiplierReg_223 = _RAND_1478[4:0];
  _RAND_1479 = {1{`RANDOM}};
  signReg_223 = _RAND_1479[0:0];
  _RAND_1480 = {1{`RANDOM}};
  multiplierReg_224 = _RAND_1480[4:0];
  _RAND_1481 = {1{`RANDOM}};
  signReg_224 = _RAND_1481[0:0];
  _RAND_1482 = {1{`RANDOM}};
  multiplierReg_225 = _RAND_1482[4:0];
  _RAND_1483 = {1{`RANDOM}};
  signReg_225 = _RAND_1483[0:0];
  _RAND_1484 = {1{`RANDOM}};
  multiplierReg_226 = _RAND_1484[4:0];
  _RAND_1485 = {1{`RANDOM}};
  signReg_226 = _RAND_1485[0:0];
  _RAND_1486 = {1{`RANDOM}};
  multiplierReg_227 = _RAND_1486[4:0];
  _RAND_1487 = {1{`RANDOM}};
  signReg_227 = _RAND_1487[0:0];
  _RAND_1488 = {1{`RANDOM}};
  multiplierReg_228 = _RAND_1488[4:0];
  _RAND_1489 = {1{`RANDOM}};
  signReg_228 = _RAND_1489[0:0];
  _RAND_1490 = {1{`RANDOM}};
  multiplierReg_229 = _RAND_1490[4:0];
  _RAND_1491 = {1{`RANDOM}};
  signReg_229 = _RAND_1491[0:0];
  _RAND_1492 = {1{`RANDOM}};
  multiplierReg_230 = _RAND_1492[4:0];
  _RAND_1493 = {1{`RANDOM}};
  signReg_230 = _RAND_1493[0:0];
  _RAND_1494 = {1{`RANDOM}};
  multiplierReg_231 = _RAND_1494[4:0];
  _RAND_1495 = {1{`RANDOM}};
  signReg_231 = _RAND_1495[0:0];
  _RAND_1496 = {1{`RANDOM}};
  multiplierReg_232 = _RAND_1496[4:0];
  _RAND_1497 = {1{`RANDOM}};
  signReg_232 = _RAND_1497[0:0];
  _RAND_1498 = {1{`RANDOM}};
  multiplierReg_233 = _RAND_1498[4:0];
  _RAND_1499 = {1{`RANDOM}};
  signReg_233 = _RAND_1499[0:0];
  _RAND_1500 = {1{`RANDOM}};
  multiplierReg_234 = _RAND_1500[4:0];
  _RAND_1501 = {1{`RANDOM}};
  signReg_234 = _RAND_1501[0:0];
  _RAND_1502 = {1{`RANDOM}};
  multiplierReg_235 = _RAND_1502[4:0];
  _RAND_1503 = {1{`RANDOM}};
  signReg_235 = _RAND_1503[0:0];
  _RAND_1504 = {1{`RANDOM}};
  multiplierReg_236 = _RAND_1504[4:0];
  _RAND_1505 = {1{`RANDOM}};
  signReg_236 = _RAND_1505[0:0];
  _RAND_1506 = {1{`RANDOM}};
  multiplierReg_237 = _RAND_1506[4:0];
  _RAND_1507 = {1{`RANDOM}};
  signReg_237 = _RAND_1507[0:0];
  _RAND_1508 = {1{`RANDOM}};
  multiplierReg_238 = _RAND_1508[4:0];
  _RAND_1509 = {1{`RANDOM}};
  signReg_238 = _RAND_1509[0:0];
  _RAND_1510 = {1{`RANDOM}};
  multiplierReg_239 = _RAND_1510[4:0];
  _RAND_1511 = {1{`RANDOM}};
  signReg_239 = _RAND_1511[0:0];
  _RAND_1512 = {1{`RANDOM}};
  multiplierReg_240 = _RAND_1512[4:0];
  _RAND_1513 = {1{`RANDOM}};
  signReg_240 = _RAND_1513[0:0];
  _RAND_1514 = {1{`RANDOM}};
  multiplierReg_241 = _RAND_1514[4:0];
  _RAND_1515 = {1{`RANDOM}};
  signReg_241 = _RAND_1515[0:0];
  _RAND_1516 = {1{`RANDOM}};
  multiplierReg_242 = _RAND_1516[4:0];
  _RAND_1517 = {1{`RANDOM}};
  signReg_242 = _RAND_1517[0:0];
  _RAND_1518 = {1{`RANDOM}};
  multiplierReg_243 = _RAND_1518[4:0];
  _RAND_1519 = {1{`RANDOM}};
  signReg_243 = _RAND_1519[0:0];
  _RAND_1520 = {1{`RANDOM}};
  multiplierReg_244 = _RAND_1520[4:0];
  _RAND_1521 = {1{`RANDOM}};
  signReg_244 = _RAND_1521[0:0];
  _RAND_1522 = {1{`RANDOM}};
  multiplierReg_245 = _RAND_1522[4:0];
  _RAND_1523 = {1{`RANDOM}};
  signReg_245 = _RAND_1523[0:0];
  _RAND_1524 = {1{`RANDOM}};
  multiplierReg_246 = _RAND_1524[4:0];
  _RAND_1525 = {1{`RANDOM}};
  signReg_246 = _RAND_1525[0:0];
  _RAND_1526 = {1{`RANDOM}};
  multiplierReg_247 = _RAND_1526[4:0];
  _RAND_1527 = {1{`RANDOM}};
  signReg_247 = _RAND_1527[0:0];
  _RAND_1528 = {1{`RANDOM}};
  multiplierReg_248 = _RAND_1528[4:0];
  _RAND_1529 = {1{`RANDOM}};
  signReg_248 = _RAND_1529[0:0];
  _RAND_1530 = {1{`RANDOM}};
  multiplierReg_249 = _RAND_1530[4:0];
  _RAND_1531 = {1{`RANDOM}};
  signReg_249 = _RAND_1531[0:0];
  _RAND_1532 = {1{`RANDOM}};
  multiplierReg_250 = _RAND_1532[4:0];
  _RAND_1533 = {1{`RANDOM}};
  signReg_250 = _RAND_1533[0:0];
  _RAND_1534 = {1{`RANDOM}};
  multiplierReg_251 = _RAND_1534[4:0];
  _RAND_1535 = {1{`RANDOM}};
  signReg_251 = _RAND_1535[0:0];
  _RAND_1536 = {1{`RANDOM}};
  multiplierReg_252 = _RAND_1536[4:0];
  _RAND_1537 = {1{`RANDOM}};
  signReg_252 = _RAND_1537[0:0];
  _RAND_1538 = {1{`RANDOM}};
  multiplierReg_253 = _RAND_1538[4:0];
  _RAND_1539 = {1{`RANDOM}};
  signReg_253 = _RAND_1539[0:0];
  _RAND_1540 = {1{`RANDOM}};
  multiplierReg_254 = _RAND_1540[4:0];
  _RAND_1541 = {1{`RANDOM}};
  signReg_254 = _RAND_1541[0:0];
  _RAND_1542 = {1{`RANDOM}};
  multiplierReg_255 = _RAND_1542[4:0];
  _RAND_1543 = {1{`RANDOM}};
  signReg_255 = _RAND_1543[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
